/****************************************************************************
 *                                                                          *
 *  FLAT VERSION of HIGH-LEVEL MODEL for c1908                              *
 *                                                                          *
 *                                                                          *
 *  Generated by: Hakan Yalcin (hyalcin@cadence.com)                        *
 *  Verified  by: Jonathan David Hauke (jhauke@eecs.umich.edu)              *
 *                                                                          *
 *                Oct 20, 1998                                              *
 *                                                                          *
****************************************************************************/
// Flat Verilog File 
module c1908g (
	in101, in104, in107, in110, in113, in116, in119, 
	in122, in125, in128, in131, in134, in137, in140, in143, 
	in146, in210, in214, in217, in221, in224, in227, in234, 
	in237, in469, in472, in475, in478, in898, in900, in902, 
	in952, in953,
	out3, out6, out9, out12, out30, out45, out48, 
	out15, out18, out21, out24, out27, out33, out36, out39, 
	out42, out75, out51, out54, out60, out63, out66, out69, 
	out72, out57);

   input
	in101, in104, in107, in110, in113, in116, in119, 
	in122, in125, in128, in131, in134, in137, in140, in143, 
	in146, in210, in214, in217, in221, in224, in227, in234, 
	in237, in469, in472, in475, in478, in898, in900, in902, 
	in952, in953;

   output
	out3, out6, out9, out12, out30, out45, out48, 
	out15, out18, out21, out24, out27, out33, out36, out39, 
	out42, out75, out51, out54, out60, out63, out66, out69, 
	out72, out57;

inv M1_UM1_0(in953, M1_Not_ContB);
inv M1_UM1_1(in237, M1_Not_ContH);
and3 M1_UM1_2(in217, in234, M1_Not_ContB, M1_temp0);
and3 M1_UM1_3(in214, M1_Not_ContH, M1_Not_ContB, M1_temp1);
and3 M1_UM1_4(in210, M1_Not_ContH, M1_Not_ContB, M1_temp2);
and2 M1_UM1_5(in227, M1_Not_ContB, M1_temp3);
and3 M1_UM1_6(in221, in234, M1_Not_ContB, M1_temp4);
and2 M1_UM1_7(in224, M1_Not_ContB, M1_temp5);
inv M1_UM1_8(in101, M1_NotInDataBus_0);
inv M1_UM1_9(in104, M1_NotInDataBus_1);
inv M1_UM1_10(in107, M1_NotInDataBus_2);
inv M1_UM1_11(in110, M1_NotInDataBus_3);
inv M1_UM1_12(in113, M1_NotInDataBus_4);
inv M1_UM1_13(in116, M1_NotInDataBus_5);
inv M1_UM1_14(in119, M1_NotInDataBus_6);
inv M1_UM1_15(in122, M1_NotInDataBus_7);
inv M1_UM1_16(in125, M1_NotInDataBus_8);
inv M1_UM1_17(in128, M1_NotInDataBus_9);
inv M1_UM1_18(in131, M1_NotInDataBus_10);
inv M1_UM1_19(in134, M1_NotInDataBus_11);
inv M1_UM1_20(in137, M1_NotInDataBus_12);
inv M1_UM1_21(in140, M1_NotInDataBus_13);
inv M1_UM1_22(in143, M1_NotInDataBus_14);
inv M1_UM1_23(in146, M1_NotInDataBus_15);
xor2 M1_UM1_46(M1_NotInDataBus_7, M1_NotInDataBus_5, M1_line46);
xor2 M1_UM1_47(M1_line46, M1_NotInDataBus_2, M1_line47);
xor2 M1_UM1_48(M1_NotInDataBus_14, M1_NotInDataBus_9, M1_line48);
xor2 M1_UM1_49(M1_line48, M1_NotInDataBus_11, M1_line49);
xor2 M1_UM1_50(M1_line47, M1_line49, M1_line50);
xor2 M1_UM1_51(M1_line50, M1_temp0, SynBits_0);
xor2 M1_UM1_38(M1_NotInDataBus_8, M1_NotInDataBus_13, M1_line38);
xor2 M1_UM1_39(M1_line38, M1_NotInDataBus_15, M1_line39);
xor2 M1_UM1_40(M1_NotInDataBus_14, M1_temp1, M1_line40);
xor2 M1_UM1_41(M1_line40, M1_NotInDataBus_10, M1_line41);
xor2 M1_UM1_42(M1_line39, M1_line41, M1_line42);
xor2 M1_UM1_43(M1_NotInDataBus_7, M1_NotInDataBus_4, M1_line43);
xor2 M1_UM1_44(M1_line43, M1_NotInDataBus_1, M1_line44);
xor2 M1_UM1_45(M1_line42, M1_line44, SynBits_1);
xor2 M1_UM1_24(M1_NotInDataBus_0, M1_temp2, M1_line24);
xor2 M1_UM1_25(M1_NotInDataBus_12, M1_NotInDataBus_11, M1_line25);
xor2 M1_UM1_26(M1_line25, M1_NotInDataBus_10, M1_line26);
inv M1_UM1_27(M1_line26, M1_line27);
xor2 M1_UM1_28(M1_NotInDataBus_15, M1_NotInDataBus_14, M1_line28);
xor2 M1_UM1_29(M1_line28, M1_NotInDataBus_9, M1_line29);
xor2 M1_UM1_30(M1_line27, M1_line29, M1_line30);
xor2 M1_UM1_31(M1_NotInDataBus_6, M1_NotInDataBus_5, M1_line31);
xor2 M1_UM1_32(M1_line31, M1_NotInDataBus_4, M1_line32);
inv M1_UM1_33(M1_line32, M1_line33);
xor2 M1_UM1_34(M1_line30, M1_line33, M1_line34);
inv M1_UM1_35(M1_line34, M1_line35);
inv M1_UM1_36(M1_line24, M1_line36);
xor2 M1_UM1_37(M1_line36, M1_line35, SynBits_2);
xor2 M1_UM1_76(M1_NotInDataBus_3, M1_NotInDataBus_13, M1_line76);
xor2 M1_UM1_77(M1_line76, M1_temp3, M1_line77);
xor2 M1_UM1_78(M1_NotInDataBus_2, M1_NotInDataBus_1, M1_line78);
xor2 M1_UM1_79(M1_line78, M1_NotInDataBus_0, M1_line79);
xor2 M1_UM1_80(M1_NotInDataBus_15, M1_NotInDataBus_14, M1_line80);
xor2 M1_UM1_81(M1_line80, M1_NotInDataBus_9, M1_line81);
inv M1_UM1_82(M1_line81, M1_line82);
xor2 M1_UM1_83(M1_line79, M1_line82, M1_line83);
xor2 M1_UM1_84(M1_line83, M1_line27, M1_line84);
inv M1_UM1_85(M1_line84, M1_line85);
xor2 M1_UM1_86(M1_line77, M1_line85, SynBits_3);
xor2 M1_UM1_52(M1_NotInDataBus_8, M1_NotInDataBus_13, M1_line52);
xor2 M1_UM1_53(M1_line52, M1_NotInDataBus_15, M1_line53);
inv M1_UM1_54(M1_line53, M1_line54);
xor2 M1_UM1_55(M1_NotInDataBus_9, M1_NotInDataBus_6, M1_line55);
xor2 M1_UM1_56(M1_line55, M1_NotInDataBus_3, M1_line56);
inv M1_UM1_57(M1_line56, M1_line57);
xor2 M1_UM1_58(M1_line54, M1_line57, M1_line58);
xor2 M1_UM1_59(M1_temp4, M1_NotInDataBus_12, M1_line59);
inv M1_UM1_60(M1_line59, M1_line60);
xor2 M1_UM1_61(M1_line58, M1_line60, SynBits_4);
xor2 M1_UM1_62(M1_line29, M1_NotInDataBus_8, M1_line62);
xor2 M1_UM1_63(M1_line62, M1_temp5, M1_line63);
inv M1_UM1_64(M1_line63, M1_line64);
xor2 M1_UM1_65(M1_NotInDataBus_2, M1_NotInDataBus_1, M1_line65);
xor2 M1_UM1_66(M1_line65, M1_NotInDataBus_0, M1_line66);
inv M1_UM1_67(M1_line66, M1_line67);
xor2 M1_UM1_68(M1_NotInDataBus_6, M1_NotInDataBus_5, M1_line68);
xor2 M1_UM1_69(M1_line68, M1_NotInDataBus_4, M1_line69);
xor2 M1_UM1_70(M1_line67, M1_line69, M1_line70);
xor2 M1_UM1_71(M1_NotInDataBus_7, M1_NotInDataBus_3, M1_line71);
inv M1_UM1_72(M1_line71, M1_line72);
xor2 M1_UM1_73(M1_line70, M1_line72, M1_line73);
xor2 M1_UM1_74(M1_line64, M1_line73, M1_line74);
inv M1_UM1_75(M1_line74, SynBits_5);
xor2 M1_UM1_87(M1_line67, M1_line69, M1_line87);
xor2 M1_UM1_88(M1_line87, M1_line72, InDBParityLo);
xor2 M1_UM1_89(M1_NotInDataBus_12, M1_NotInDataBus_11, M1_line89);
xor2 M1_UM1_90(M1_line89, M1_NotInDataBus_10, M1_line90);
xor2 M1_UM1_91(M1_line82, M1_line90, M1_line91);
xor2 M1_UM1_92(M1_NotInDataBus_13, M1_NotInDataBus_8, M1_line92);
inv M1_UM1_93(M1_line92, M1_line93);
xor2 M1_UM1_94(M1_line91, M1_line93, InDBParityHi);
inv M2_UM2_0(in902, M2_Not_ContE);
and2 M2_UM2_1(SynBits_0, M2_Not_ContE, M2_temp0);
and2 M2_UM2_2(SynBits_1, M2_Not_ContE, M2_temp1);
and2 M2_UM2_3(SynBits_2, M2_Not_ContE, M2_temp2);
and2 M2_UM2_4(SynBits_3, M2_Not_ContE, M2_temp3);
and2 M2_UM2_5(SynBits_4, M2_Not_ContE, M2_temp4);
and2 M2_UM2_6(SynBits_5, M2_Not_ContE, M2_temp5);
nand2 M2_UM2_7(in234, M2_Not_ContE, M2_line7);
and2 M2_UM2_8(in217, M2_line7, AllExtSynBits_4);
inv M2_UM2_9(in237, M2_Not_ContH);
nand2 M2_UM2_10(M2_Not_ContH, M2_Not_ContE, M2_line10);
and2 M2_UM2_11(M2_line10, in210, AllExtSynBits_5);
nand2 M2_UM2_12(in214, M2_line10, ContIntM);
nand2 M2_UM2_13(in221, M2_line7, ContIntP);
xor2 M2_UM2_14(M2_temp0, in478, NewSynBits_0);
xor2 M2_UM2_15(M2_temp1, in475, NewSynBits_1);
xor2 M2_UM2_16(M2_temp2, in472, NewSynBits_2);
xor2 M2_UM2_17(M2_temp3, in469, NewSynBits_3);
xor2 M2_UM2_18(M2_temp4, AllExtSynBits_4, NewSynBits_4);
xor2 M2_UM2_19(M2_temp5, AllExtSynBits_5, NewSynBits_5);
inv M2_UM2_20(NewSynBits_0, Not_NewSynBits_0);
inv M2_UM2_21(NewSynBits_1, Not_NewSynBits_1);
inv M2_UM2_22(NewSynBits_2, Not_NewSynBits_2);
inv M2_UM2_23(NewSynBits_3, Not_NewSynBits_3);
inv M2_UM2_24(NewSynBits_4, Not_NewSynBits_4);
inv M2_UM2_25(NewSynBits_5, Not_NewSynBits_5);
inv M3_UM3_0(in898, M3_Not_ContK);
inv M3_UM3_1(in900, M3_Not_ContL);
inv M3_UM3_2(in953, M3_Not_ContB);
nand2 M3_UM3_3(in234, in237, M3_NotGH);
nand4 M3_UM3_4(M3_Not_ContK, in902, in953, M3_NotGH, M3_line4);
nand3 M3_UM3_5(in952, M3_Not_ContB, M3_NotGH, M3_line5);
nand2 M3_UM3_6(M3_line4, M3_line5, M3_ContIntLo);
nand4 M3_UM3_7(M3_Not_ContL, in902, in953, M3_NotGH, M3_line7);
nand2 M3_UM3_8(M3_line7, M3_line5, M3_ContIntHi);
and2 M3_UM3_9(ContIntM, NewSynBits_5, ProductSyn_0);
and2 M3_UM3_10(Not_NewSynBits_0, Not_NewSynBits_1, ProductSyn_1);
and2 M3_UM3_11(Not_NewSynBits_4, Not_NewSynBits_2, ProductSyn_2);
and2 M3_UM3_12(Not_NewSynBits_0, NewSynBits_1, ProductSyn_3);
and2 M3_UM3_13(NewSynBits_0, Not_NewSynBits_1, ProductSyn_4);
and2 M3_UM3_14(NewSynBits_4, Not_NewSynBits_2, ProductSyn_5);
and2 M3_UM3_15(ContIntP, Not_NewSynBits_3, ProductSyn_6);
and2 M3_UM3_16(NewSynBits_4, NewSynBits_2, ProductSyn_7);
and2 M3_UM3_17(ContIntM, Not_NewSynBits_5, ProductSyn_8);
and2 M3_UM3_18(Not_NewSynBits_4, NewSynBits_2, ProductSyn_9);
and2 M3_UM3_19(ContIntP, NewSynBits_3, ProductSyn_10);
and2 M3_UM3_20(NewSynBits_0, NewSynBits_1, ProductSyn_11);
and5 M3_UM3_21(ProductSyn_0, ProductSyn_10, ProductSyn_9, ProductSyn_1, M3_ContIntLo, DecodedSyn_0);
and5 M3_UM3_22(ProductSyn_0, ProductSyn_10, ProductSyn_2, ProductSyn_3, M3_ContIntLo, DecodedSyn_1);
and5 M3_UM3_23(ProductSyn_0, ProductSyn_10, ProductSyn_2, ProductSyn_4, M3_ContIntLo, DecodedSyn_2);
and5 M3_UM3_24(ProductSyn_0, ProductSyn_10, ProductSyn_5, ProductSyn_1, M3_ContIntLo, DecodedSyn_3);
and5 M3_UM3_25(ProductSyn_0, ProductSyn_6, ProductSyn_9, ProductSyn_3, M3_ContIntLo, DecodedSyn_4);
and5 M3_UM3_26(ProductSyn_0, ProductSyn_6, ProductSyn_9, ProductSyn_4, M3_ContIntLo, DecodedSyn_5);
and5 M3_UM3_27(ProductSyn_0, ProductSyn_6, ProductSyn_7, ProductSyn_1, M3_ContIntLo, DecodedSyn_6);
and5 M3_UM3_28(ProductSyn_0, ProductSyn_6, ProductSyn_2, ProductSyn_11, M3_ContIntLo, DecodedSyn_7);
and5 M3_UM3_29(ProductSyn_0, ProductSyn_6, ProductSyn_5, ProductSyn_3, M3_ContIntHi, DecodedSyn_8);
and5 M3_UM3_30(ProductSyn_0, ProductSyn_10, ProductSyn_7, ProductSyn_4, M3_ContIntHi, DecodedSyn_9);
and5 M3_UM3_31(ProductSyn_8, ProductSyn_10, ProductSyn_9, ProductSyn_3, M3_ContIntHi, DecodedSyn_10);
and5 M3_UM3_32(ProductSyn_8, ProductSyn_10, ProductSyn_9, ProductSyn_4, M3_ContIntHi, DecodedSyn_11);
and5 M3_UM3_33(ProductSyn_8, ProductSyn_10, ProductSyn_7, ProductSyn_1, M3_ContIntHi, DecodedSyn_12);
and5 M3_UM3_34(ProductSyn_8, ProductSyn_10, ProductSyn_5, ProductSyn_3, M3_ContIntHi, DecodedSyn_13);
and5 M3_UM3_35(ProductSyn_0, ProductSyn_10, ProductSyn_9, ProductSyn_11, M3_ContIntHi, DecodedSyn_14);
and5 M3_UM3_36(ProductSyn_0, ProductSyn_10, ProductSyn_7, ProductSyn_3, M3_ContIntHi, DecodedSyn_15);
or8 M3_UM3_37(DecodedSyn_0, DecodedSyn_1, DecodedSyn_2, DecodedSyn_3, DecodedSyn_4, DecodedSyn_5, DecodedSyn_6, DecodedSyn_7, CorrectionFlagLo);
or8 M3_UM3_38(DecodedSyn_8, DecodedSyn_9, DecodedSyn_10, DecodedSyn_11, DecodedSyn_12, DecodedSyn_13, DecodedSyn_14, DecodedSyn_15, CorrectionFlagHi);
or2 M3_UM3_39(CorrectionFlagLo, CorrectionFlagHi, CorrectionFlag);
xor2 M4_UM4_0(in101, DecodedSyn_0, out3);
xor2 M4_UM4_1(in104, DecodedSyn_1, out6);
xor2 M4_UM4_2(in107, DecodedSyn_2, out9);
xor2 M4_UM4_3(in110, DecodedSyn_3, out12);
xor2 M4_UM4_4(in113, DecodedSyn_4, out15);
xor2 M4_UM4_5(in116, DecodedSyn_5, out18);
xor2 M4_UM4_6(in119, DecodedSyn_6, out21);
xor2 M4_UM4_7(in122, DecodedSyn_7, out24);
xor2 M4_UM4_8(in125, DecodedSyn_8, out27);
xor2 M4_UM4_9(in128, DecodedSyn_9, out30);
xor2 M4_UM4_10(in131, DecodedSyn_10, out33);
xor2 M4_UM4_11(in134, DecodedSyn_11, out36);
xor2 M4_UM4_12(in137, DecodedSyn_12, out39);
xor2 M4_UM4_13(in140, DecodedSyn_13, out42);
xor2 M4_UM4_14(in143, DecodedSyn_14, out45);
xor2 M4_UM4_15(in146, DecodedSyn_15, out48);
inv M5_UM5_0(in952, M5_Not_ContF);
and3 M5_UM5_1_SCS_0(in478, in902, CorrectionFlag, M5_UM5_1_line0);
xor2 M5_UM5_1_SCS_1(SynBits_0, M5_UM5_1_line0, M5_UM5_1_line1);
nand2 M5_UM5_1_SCS_2(M5_Not_ContF, in953, M5_UM5_1_line2);
and2 M5_UM5_1_SCS_3(M5_UM5_1_line2, M5_UM5_1_line1, out63);
and3 M5_UM5_2_SCS_0(in475, in902, CorrectionFlag, M5_UM5_2_line0);
xor2 M5_UM5_2_SCS_1(SynBits_1, M5_UM5_2_line0, M5_UM5_2_line1);
nand2 M5_UM5_2_SCS_2(M5_Not_ContF, in953, M5_UM5_2_line2);
and2 M5_UM5_2_SCS_3(M5_UM5_2_line2, M5_UM5_2_line1, out60);
and3 M5_UM5_3_SCS_0(in472, in902, CorrectionFlag, M5_UM5_3_line0);
xor2 M5_UM5_3_SCS_1(SynBits_2, M5_UM5_3_line0, M5_UM5_3_line1);
nand2 M5_UM5_3_SCS_2(M5_Not_ContF, in953, M5_UM5_3_line2);
and2 M5_UM5_3_SCS_3(M5_UM5_3_line2, M5_UM5_3_line1, out57);
and3 M5_UM5_4_SCS_0(in469, in902, CorrectionFlag, M5_UM5_4_line0);
xor2 M5_UM5_4_SCS_1(SynBits_3, M5_UM5_4_line0, M5_UM5_4_line1);
nand2 M5_UM5_4_SCS_2(M5_Not_ContF, in953, M5_UM5_4_line2);
and2 M5_UM5_4_SCS_3(M5_UM5_4_line2, M5_UM5_4_line1, out54);
and3 M5_UM5_5_SCS_0(AllExtSynBits_4, in902, CorrectionFlag, M5_UM5_5_line0);
xor2 M5_UM5_5_SCS_1(SynBits_4, M5_UM5_5_line0, M5_UM5_5_line1);
nand2 M5_UM5_5_SCS_2(M5_Not_ContF, in953, M5_UM5_5_line2);
and2 M5_UM5_5_SCS_3(M5_UM5_5_line2, M5_UM5_5_line1, out66);
and3 M5_UM5_6_SCS_0(AllExtSynBits_5, in902, CorrectionFlag, M5_UM5_6_line0);
xor2 M5_UM5_6_SCS_1(SynBits_5, M5_UM5_6_line0, M5_UM5_6_line1);
nand2 M5_UM5_6_SCS_2(M5_Not_ContF, in953, M5_UM5_6_line2);
and2 M5_UM5_6_SCS_3(M5_UM5_6_line2, M5_UM5_6_line1, out51);
inv M6_UM6_7_0(in953, M6_Not_ContB);
inv M6_UM6_7_1(in900, M6_Not_Cont_N);
inv M6_UM6_7_2(InDBParityHi, M6_Not_InDBParity_N);
nand2 M6_UM6_7_3(in953, M6_Not_Cont_N, M6_line3);
and2 M6_UM6_7_4(M6_line3, M6_Not_InDBParity_N, M6_line4);
and2 M6_UM6_7_5(CorrectionFlagHi, M6_Not_ContB, M6_line5);
xor2 M6_UM6_7_6(M6_line5, M6_line4, M6_line6);
nand2 M6_UM6_7_7(in227, in900, M6_line7);
and2 M6_UM6_7_8(M6_line7, in953, M6_line8);
xor2 M6_UM6_7_9(M6_line6, M6_line8, out72);
inv M7_UM6_7_0(in953, M7_Not_ContB);
inv M7_UM6_7_1(in898, M7_Not_Cont_N);
inv M7_UM6_7_2(InDBParityLo, M7_Not_InDBParity_N);
nand2 M7_UM6_7_3(in953, M7_Not_Cont_N, M7_line3);
and2 M7_UM6_7_4(M7_line3, M7_Not_InDBParity_N, M7_line4);
and2 M7_UM6_7_5(CorrectionFlagLo, M7_Not_ContB, M7_line5);
xor2 M7_UM6_7_6(M7_line5, M7_line4, M7_line6);
nand2 M7_UM6_7_7(in224, in898, M7_line7);
and2 M7_UM6_7_8(M7_line7, in953, M7_line8);
xor2 M7_UM6_7_9(M7_line6, M7_line8, out69);
inv M8_UM8_0(in237, M8_Not_ContH);
inv M8_UM8_1(in902, M8_Not_ContE);
inv M8_UM8_2(in953, M8_Not_ContB);
inv M8_UM8_3(in952, M8_Not_ContF);
inv M8_UM8_4(ContIntM, M8_NotM);
inv M8_UM8_5(ContIntP, M8_NotP);
nand2 M8_UM8_6(in234, in237, M8_NotGH);
and3 M8_UM8_7(in952, M8_Not_ContB, M8_NotGH, M8_ContIntUE);
and2 M8_UM8_8_UEG_0(M8_NotP, Not_NewSynBits_3, M8_UM8_8_line0);
and2 M8_UM8_8_UEG_1(M8_NotM, Not_NewSynBits_5, M8_UM8_8_line1);
nand5 M8_UM8_8_UEG_2(ProductSyn_0, ProductSyn_6, ProductSyn_2, ProductSyn_1, M8_ContIntUE, M8_UM8_8_line2);
nand5 M8_UM8_8_UEG_3(ProductSyn_8, ProductSyn_10, ProductSyn_2, ProductSyn_1, M8_ContIntUE, M8_UM8_8_line3);
nand5 M8_UM8_8_UEG_4(ProductSyn_8, ProductSyn_6, ProductSyn_9, ProductSyn_1, M8_ContIntUE, M8_UM8_8_line4);
nand5 M8_UM8_8_UEG_5(ProductSyn_8, ProductSyn_6, ProductSyn_2, ProductSyn_3, M8_ContIntUE, M8_UM8_8_line5);
nand5 M8_UM8_8_UEG_6(ProductSyn_8, ProductSyn_6, ProductSyn_2, ProductSyn_4, M8_ContIntUE, M8_UM8_8_line6);
nand5 M8_UM8_8_UEG_7(ProductSyn_8, ProductSyn_6, ProductSyn_5, ProductSyn_1, M8_ContIntUE, M8_UM8_8_line7);
nand5 M8_UM8_8_UEG_8(ProductSyn_8, M8_UM8_8_line0, ProductSyn_2, ProductSyn_1, M8_ContIntUE, M8_UM8_8_line8);
nand5 M8_UM8_8_UEG_9(M8_UM8_8_line1, ProductSyn_6, ProductSyn_2, ProductSyn_1, M8_ContIntUE, M8_UM8_8_line9);
and8 M8_UM8_8_UEG_10(M8_UM8_8_line2, M8_UM8_8_line3, M8_UM8_8_line4, M8_UM8_8_line5, M8_UM8_8_line6, M8_UM8_8_line7, M8_UM8_8_line8, M8_UM8_8_line9, M8_UESignal);
nand2 M8_UM8_9(M8_Not_ContH, M8_Not_ContE, M8_line9);
nand2 M8_UM8_10(in214, M8_line9, M8_line10);
nand2 M8_UM8_11(in234, M8_Not_ContE, M8_line11);
nand2 M8_UM8_12(in221, M8_line11, M8_line12);
nand8 M8_UM8_13(Not_NewSynBits_0, Not_NewSynBits_1, Not_NewSynBits_2, Not_NewSynBits_3, Not_NewSynBits_4, Not_NewSynBits_5, M8_line10, M8_line12, M8_ErrorFREE);
inv M8_UM8_14(CorrectionFlagHi, M8_NotCorrFlagHi);
inv M8_UM8_15(CorrectionFlagLo, M8_NotCorrFlagLo);
and3 M8_UM8_16(M8_NotCorrFlagLo, M8_NotCorrFlagHi, M8_UESignal, M8_line16);
and4 M8_UM8_17(M8_Not_ContB, M8_ErrorFREE, in952, M8_line16, M8_line17);
and3 M8_UM8_18(M8_Not_ContB, M8_ErrorFREE, M8_Not_ContF, M8_line18);
nor2 M8_UM8_19(M8_line18, M8_line17, out75);


endmodule