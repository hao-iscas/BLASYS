module dec_tb;
reg [7:0] pi;
wire [255:0] po;
dec dut( pi[0], pi[1], pi[2], pi[3], pi[4], pi[5], pi[6], pi[7], po[0], po[1], po[2], po[3], po[4], po[5], po[6], po[7], po[8], po[9], po[10], po[11], po[12], po[13], po[14], po[15], po[16], po[17], po[18], po[19], po[20], po[21], po[22], po[23], po[24], po[25], po[26], po[27], po[28], po[29], po[30], po[31], po[32], po[33], po[34], po[35], po[36], po[37], po[38], po[39], po[40], po[41], po[42], po[43], po[44], po[45], po[46], po[47], po[48], po[49], po[50], po[51], po[52], po[53], po[54], po[55], po[56], po[57], po[58], po[59], po[60], po[61], po[62], po[63], po[64], po[65], po[66], po[67], po[68], po[69], po[70], po[71], po[72], po[73], po[74], po[75], po[76], po[77], po[78], po[79], po[80], po[81], po[82], po[83], po[84], po[85], po[86], po[87], po[88], po[89], po[90], po[91], po[92], po[93], po[94], po[95], po[96], po[97], po[98], po[99], po[100], po[101], po[102], po[103], po[104], po[105], po[106], po[107], po[108], po[109], po[110], po[111], po[112], po[113], po[114], po[115], po[116], po[117], po[118], po[119], po[120], po[121], po[122], po[123], po[124], po[125], po[126], po[127], po[128], po[129], po[130], po[131], po[132], po[133], po[134], po[135], po[136], po[137], po[138], po[139], po[140], po[141], po[142], po[143], po[144], po[145], po[146], po[147], po[148], po[149], po[150], po[151], po[152], po[153], po[154], po[155], po[156], po[157], po[158], po[159], po[160], po[161], po[162], po[163], po[164], po[165], po[166], po[167], po[168], po[169], po[170], po[171], po[172], po[173], po[174], po[175], po[176], po[177], po[178], po[179], po[180], po[181], po[182], po[183], po[184], po[185], po[186], po[187], po[188], po[189], po[190], po[191], po[192], po[193], po[194], po[195], po[196], po[197], po[198], po[199], po[200], po[201], po[202], po[203], po[204], po[205], po[206], po[207], po[208], po[209], po[210], po[211], po[212], po[213], po[214], po[215], po[216], po[217], po[218], po[219], po[220], po[221], po[222], po[223], po[224], po[225], po[226], po[227], po[228], po[229], po[230], po[231], po[232], po[233], po[234], po[235], po[236], po[237], po[238], po[239], po[240], po[241], po[242], po[243], po[244], po[245], po[246], po[247], po[248], po[249], po[250], po[251], po[252], po[253], po[254], po[255]);
initial
begin
#1 pi=8'b00000000;
#1 $display("%b", po);
#1 pi=8'b00000001;
#1 $display("%b", po);
#1 pi=8'b00000010;
#1 $display("%b", po);
#1 pi=8'b00000011;
#1 $display("%b", po);
#1 pi=8'b00000100;
#1 $display("%b", po);
#1 pi=8'b00000101;
#1 $display("%b", po);
#1 pi=8'b00000110;
#1 $display("%b", po);
#1 pi=8'b00000111;
#1 $display("%b", po);
#1 pi=8'b00001000;
#1 $display("%b", po);
#1 pi=8'b00001001;
#1 $display("%b", po);
#1 pi=8'b00001010;
#1 $display("%b", po);
#1 pi=8'b00001011;
#1 $display("%b", po);
#1 pi=8'b00001100;
#1 $display("%b", po);
#1 pi=8'b00001101;
#1 $display("%b", po);
#1 pi=8'b00001110;
#1 $display("%b", po);
#1 pi=8'b00001111;
#1 $display("%b", po);
#1 pi=8'b00010000;
#1 $display("%b", po);
#1 pi=8'b00010001;
#1 $display("%b", po);
#1 pi=8'b00010010;
#1 $display("%b", po);
#1 pi=8'b00010011;
#1 $display("%b", po);
#1 pi=8'b00010100;
#1 $display("%b", po);
#1 pi=8'b00010101;
#1 $display("%b", po);
#1 pi=8'b00010110;
#1 $display("%b", po);
#1 pi=8'b00010111;
#1 $display("%b", po);
#1 pi=8'b00011000;
#1 $display("%b", po);
#1 pi=8'b00011001;
#1 $display("%b", po);
#1 pi=8'b00011010;
#1 $display("%b", po);
#1 pi=8'b00011011;
#1 $display("%b", po);
#1 pi=8'b00011100;
#1 $display("%b", po);
#1 pi=8'b00011101;
#1 $display("%b", po);
#1 pi=8'b00011110;
#1 $display("%b", po);
#1 pi=8'b00011111;
#1 $display("%b", po);
#1 pi=8'b00100000;
#1 $display("%b", po);
#1 pi=8'b00100001;
#1 $display("%b", po);
#1 pi=8'b00100010;
#1 $display("%b", po);
#1 pi=8'b00100011;
#1 $display("%b", po);
#1 pi=8'b00100100;
#1 $display("%b", po);
#1 pi=8'b00100101;
#1 $display("%b", po);
#1 pi=8'b00100110;
#1 $display("%b", po);
#1 pi=8'b00100111;
#1 $display("%b", po);
#1 pi=8'b00101000;
#1 $display("%b", po);
#1 pi=8'b00101001;
#1 $display("%b", po);
#1 pi=8'b00101010;
#1 $display("%b", po);
#1 pi=8'b00101011;
#1 $display("%b", po);
#1 pi=8'b00101100;
#1 $display("%b", po);
#1 pi=8'b00101101;
#1 $display("%b", po);
#1 pi=8'b00101110;
#1 $display("%b", po);
#1 pi=8'b00101111;
#1 $display("%b", po);
#1 pi=8'b00110000;
#1 $display("%b", po);
#1 pi=8'b00110001;
#1 $display("%b", po);
#1 pi=8'b00110010;
#1 $display("%b", po);
#1 pi=8'b00110011;
#1 $display("%b", po);
#1 pi=8'b00110100;
#1 $display("%b", po);
#1 pi=8'b00110101;
#1 $display("%b", po);
#1 pi=8'b00110110;
#1 $display("%b", po);
#1 pi=8'b00110111;
#1 $display("%b", po);
#1 pi=8'b00111000;
#1 $display("%b", po);
#1 pi=8'b00111001;
#1 $display("%b", po);
#1 pi=8'b00111010;
#1 $display("%b", po);
#1 pi=8'b00111011;
#1 $display("%b", po);
#1 pi=8'b00111100;
#1 $display("%b", po);
#1 pi=8'b00111101;
#1 $display("%b", po);
#1 pi=8'b00111110;
#1 $display("%b", po);
#1 pi=8'b00111111;
#1 $display("%b", po);
#1 pi=8'b01000000;
#1 $display("%b", po);
#1 pi=8'b01000001;
#1 $display("%b", po);
#1 pi=8'b01000010;
#1 $display("%b", po);
#1 pi=8'b01000011;
#1 $display("%b", po);
#1 pi=8'b01000100;
#1 $display("%b", po);
#1 pi=8'b01000101;
#1 $display("%b", po);
#1 pi=8'b01000110;
#1 $display("%b", po);
#1 pi=8'b01000111;
#1 $display("%b", po);
#1 pi=8'b01001000;
#1 $display("%b", po);
#1 pi=8'b01001001;
#1 $display("%b", po);
#1 pi=8'b01001010;
#1 $display("%b", po);
#1 pi=8'b01001011;
#1 $display("%b", po);
#1 pi=8'b01001100;
#1 $display("%b", po);
#1 pi=8'b01001101;
#1 $display("%b", po);
#1 pi=8'b01001110;
#1 $display("%b", po);
#1 pi=8'b01001111;
#1 $display("%b", po);
#1 pi=8'b01010000;
#1 $display("%b", po);
#1 pi=8'b01010001;
#1 $display("%b", po);
#1 pi=8'b01010010;
#1 $display("%b", po);
#1 pi=8'b01010011;
#1 $display("%b", po);
#1 pi=8'b01010100;
#1 $display("%b", po);
#1 pi=8'b01010101;
#1 $display("%b", po);
#1 pi=8'b01010110;
#1 $display("%b", po);
#1 pi=8'b01010111;
#1 $display("%b", po);
#1 pi=8'b01011000;
#1 $display("%b", po);
#1 pi=8'b01011001;
#1 $display("%b", po);
#1 pi=8'b01011010;
#1 $display("%b", po);
#1 pi=8'b01011011;
#1 $display("%b", po);
#1 pi=8'b01011100;
#1 $display("%b", po);
#1 pi=8'b01011101;
#1 $display("%b", po);
#1 pi=8'b01011110;
#1 $display("%b", po);
#1 pi=8'b01011111;
#1 $display("%b", po);
#1 pi=8'b01100000;
#1 $display("%b", po);
#1 pi=8'b01100001;
#1 $display("%b", po);
#1 pi=8'b01100010;
#1 $display("%b", po);
#1 pi=8'b01100011;
#1 $display("%b", po);
#1 pi=8'b01100100;
#1 $display("%b", po);
#1 pi=8'b01100101;
#1 $display("%b", po);
#1 pi=8'b01100110;
#1 $display("%b", po);
#1 pi=8'b01100111;
#1 $display("%b", po);
#1 pi=8'b01101000;
#1 $display("%b", po);
#1 pi=8'b01101001;
#1 $display("%b", po);
#1 pi=8'b01101010;
#1 $display("%b", po);
#1 pi=8'b01101011;
#1 $display("%b", po);
#1 pi=8'b01101100;
#1 $display("%b", po);
#1 pi=8'b01101101;
#1 $display("%b", po);
#1 pi=8'b01101110;
#1 $display("%b", po);
#1 pi=8'b01101111;
#1 $display("%b", po);
#1 pi=8'b01110000;
#1 $display("%b", po);
#1 pi=8'b01110001;
#1 $display("%b", po);
#1 pi=8'b01110010;
#1 $display("%b", po);
#1 pi=8'b01110011;
#1 $display("%b", po);
#1 pi=8'b01110100;
#1 $display("%b", po);
#1 pi=8'b01110101;
#1 $display("%b", po);
#1 pi=8'b01110110;
#1 $display("%b", po);
#1 pi=8'b01110111;
#1 $display("%b", po);
#1 pi=8'b01111000;
#1 $display("%b", po);
#1 pi=8'b01111001;
#1 $display("%b", po);
#1 pi=8'b01111010;
#1 $display("%b", po);
#1 pi=8'b01111011;
#1 $display("%b", po);
#1 pi=8'b01111100;
#1 $display("%b", po);
#1 pi=8'b01111101;
#1 $display("%b", po);
#1 pi=8'b01111110;
#1 $display("%b", po);
#1 pi=8'b01111111;
#1 $display("%b", po);
#1 pi=8'b10000000;
#1 $display("%b", po);
#1 pi=8'b10000001;
#1 $display("%b", po);
#1 pi=8'b10000010;
#1 $display("%b", po);
#1 pi=8'b10000011;
#1 $display("%b", po);
#1 pi=8'b10000100;
#1 $display("%b", po);
#1 pi=8'b10000101;
#1 $display("%b", po);
#1 pi=8'b10000110;
#1 $display("%b", po);
#1 pi=8'b10000111;
#1 $display("%b", po);
#1 pi=8'b10001000;
#1 $display("%b", po);
#1 pi=8'b10001001;
#1 $display("%b", po);
#1 pi=8'b10001010;
#1 $display("%b", po);
#1 pi=8'b10001011;
#1 $display("%b", po);
#1 pi=8'b10001100;
#1 $display("%b", po);
#1 pi=8'b10001101;
#1 $display("%b", po);
#1 pi=8'b10001110;
#1 $display("%b", po);
#1 pi=8'b10001111;
#1 $display("%b", po);
#1 pi=8'b10010000;
#1 $display("%b", po);
#1 pi=8'b10010001;
#1 $display("%b", po);
#1 pi=8'b10010010;
#1 $display("%b", po);
#1 pi=8'b10010011;
#1 $display("%b", po);
#1 pi=8'b10010100;
#1 $display("%b", po);
#1 pi=8'b10010101;
#1 $display("%b", po);
#1 pi=8'b10010110;
#1 $display("%b", po);
#1 pi=8'b10010111;
#1 $display("%b", po);
#1 pi=8'b10011000;
#1 $display("%b", po);
#1 pi=8'b10011001;
#1 $display("%b", po);
#1 pi=8'b10011010;
#1 $display("%b", po);
#1 pi=8'b10011011;
#1 $display("%b", po);
#1 pi=8'b10011100;
#1 $display("%b", po);
#1 pi=8'b10011101;
#1 $display("%b", po);
#1 pi=8'b10011110;
#1 $display("%b", po);
#1 pi=8'b10011111;
#1 $display("%b", po);
#1 pi=8'b10100000;
#1 $display("%b", po);
#1 pi=8'b10100001;
#1 $display("%b", po);
#1 pi=8'b10100010;
#1 $display("%b", po);
#1 pi=8'b10100011;
#1 $display("%b", po);
#1 pi=8'b10100100;
#1 $display("%b", po);
#1 pi=8'b10100101;
#1 $display("%b", po);
#1 pi=8'b10100110;
#1 $display("%b", po);
#1 pi=8'b10100111;
#1 $display("%b", po);
#1 pi=8'b10101000;
#1 $display("%b", po);
#1 pi=8'b10101001;
#1 $display("%b", po);
#1 pi=8'b10101010;
#1 $display("%b", po);
#1 pi=8'b10101011;
#1 $display("%b", po);
#1 pi=8'b10101100;
#1 $display("%b", po);
#1 pi=8'b10101101;
#1 $display("%b", po);
#1 pi=8'b10101110;
#1 $display("%b", po);
#1 pi=8'b10101111;
#1 $display("%b", po);
#1 pi=8'b10110000;
#1 $display("%b", po);
#1 pi=8'b10110001;
#1 $display("%b", po);
#1 pi=8'b10110010;
#1 $display("%b", po);
#1 pi=8'b10110011;
#1 $display("%b", po);
#1 pi=8'b10110100;
#1 $display("%b", po);
#1 pi=8'b10110101;
#1 $display("%b", po);
#1 pi=8'b10110110;
#1 $display("%b", po);
#1 pi=8'b10110111;
#1 $display("%b", po);
#1 pi=8'b10111000;
#1 $display("%b", po);
#1 pi=8'b10111001;
#1 $display("%b", po);
#1 pi=8'b10111010;
#1 $display("%b", po);
#1 pi=8'b10111011;
#1 $display("%b", po);
#1 pi=8'b10111100;
#1 $display("%b", po);
#1 pi=8'b10111101;
#1 $display("%b", po);
#1 pi=8'b10111110;
#1 $display("%b", po);
#1 pi=8'b10111111;
#1 $display("%b", po);
#1 pi=8'b11000000;
#1 $display("%b", po);
#1 pi=8'b11000001;
#1 $display("%b", po);
#1 pi=8'b11000010;
#1 $display("%b", po);
#1 pi=8'b11000011;
#1 $display("%b", po);
#1 pi=8'b11000100;
#1 $display("%b", po);
#1 pi=8'b11000101;
#1 $display("%b", po);
#1 pi=8'b11000110;
#1 $display("%b", po);
#1 pi=8'b11000111;
#1 $display("%b", po);
#1 pi=8'b11001000;
#1 $display("%b", po);
#1 pi=8'b11001001;
#1 $display("%b", po);
#1 pi=8'b11001010;
#1 $display("%b", po);
#1 pi=8'b11001011;
#1 $display("%b", po);
#1 pi=8'b11001100;
#1 $display("%b", po);
#1 pi=8'b11001101;
#1 $display("%b", po);
#1 pi=8'b11001110;
#1 $display("%b", po);
#1 pi=8'b11001111;
#1 $display("%b", po);
#1 pi=8'b11010000;
#1 $display("%b", po);
#1 pi=8'b11010001;
#1 $display("%b", po);
#1 pi=8'b11010010;
#1 $display("%b", po);
#1 pi=8'b11010011;
#1 $display("%b", po);
#1 pi=8'b11010100;
#1 $display("%b", po);
#1 pi=8'b11010101;
#1 $display("%b", po);
#1 pi=8'b11010110;
#1 $display("%b", po);
#1 pi=8'b11010111;
#1 $display("%b", po);
#1 pi=8'b11011000;
#1 $display("%b", po);
#1 pi=8'b11011001;
#1 $display("%b", po);
#1 pi=8'b11011010;
#1 $display("%b", po);
#1 pi=8'b11011011;
#1 $display("%b", po);
#1 pi=8'b11011100;
#1 $display("%b", po);
#1 pi=8'b11011101;
#1 $display("%b", po);
#1 pi=8'b11011110;
#1 $display("%b", po);
#1 pi=8'b11011111;
#1 $display("%b", po);
#1 pi=8'b11100000;
#1 $display("%b", po);
#1 pi=8'b11100001;
#1 $display("%b", po);
#1 pi=8'b11100010;
#1 $display("%b", po);
#1 pi=8'b11100011;
#1 $display("%b", po);
#1 pi=8'b11100100;
#1 $display("%b", po);
#1 pi=8'b11100101;
#1 $display("%b", po);
#1 pi=8'b11100110;
#1 $display("%b", po);
#1 pi=8'b11100111;
#1 $display("%b", po);
#1 pi=8'b11101000;
#1 $display("%b", po);
#1 pi=8'b11101001;
#1 $display("%b", po);
#1 pi=8'b11101010;
#1 $display("%b", po);
#1 pi=8'b11101011;
#1 $display("%b", po);
#1 pi=8'b11101100;
#1 $display("%b", po);
#1 pi=8'b11101101;
#1 $display("%b", po);
#1 pi=8'b11101110;
#1 $display("%b", po);
#1 pi=8'b11101111;
#1 $display("%b", po);
#1 pi=8'b11110000;
#1 $display("%b", po);
#1 pi=8'b11110001;
#1 $display("%b", po);
#1 pi=8'b11110010;
#1 $display("%b", po);
#1 pi=8'b11110011;
#1 $display("%b", po);
#1 pi=8'b11110100;
#1 $display("%b", po);
#1 pi=8'b11110101;
#1 $display("%b", po);
#1 pi=8'b11110110;
#1 $display("%b", po);
#1 pi=8'b11110111;
#1 $display("%b", po);
#1 pi=8'b11111000;
#1 $display("%b", po);
#1 pi=8'b11111001;
#1 $display("%b", po);
#1 pi=8'b11111010;
#1 $display("%b", po);
#1 pi=8'b11111011;
#1 $display("%b", po);
#1 pi=8'b11111100;
#1 $display("%b", po);
#1 pi=8'b11111101;
#1 $display("%b", po);
#1 pi=8'b11111110;
#1 $display("%b", po);
#1 pi=8'b11111111;
#1 $display("%b", po);
end
endmodule
