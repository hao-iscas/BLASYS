/****************************************************************************
 *                                                                          *
 *  FLAT VERSION of HIGH-LEVEL MODEL for c5315                              *
 *                                                                          *
 *                                                                          *
 *  Generated by: Hakan Yalcin (hyalcin@cadence.com)                        *
 *  Verified  by: Jonathan David Hauke (jhauke@eecs.umich.edu)              *
 *                                                                          *
 *                Oct 20, 1998                                              *
 *                                                                          *
****************************************************************************/

// Flat Verilog File 
module c5315g (
	in293, in302, in308, in316, in324, in341, in351, 
	in361, in299, in307, in315, in323, in331, in338, in348, 
	in358, in366, in206, in210, in218, in226, in234, in257, 
	in265, in273, in281, in209, in217, in225, in233, in241, 
	in264, in272, in280, in288, in54, in4, in2174, in1497, 
	in332, in335, in479, in490, in503, in514, in523, in534, 
	in446, in457, in468, in422, in435, in389, in400, in411, 
	in374, in191, in200, in194, in197, in203, in149, in155, 
	in188, in182, in161, in170, in164, in167, in173, in146, 
	in152, in158, in185, in109, in43, in46, in100, in91, 
	in76, in73, in67, in11, in106, in37, in49, in103, 
	in40, in20, in17, in70, in61, in123, in52, in121, 
	in116, in112, in130, in119, in129, in131, in115, in122, 
	in114, in53, in113, in128, in127, in126, in117, in176, 
	in179, in14, in64, in248, in251, in242, in254, in3552, 
	in3550, in3546, in3548, in120, in94, in118, in97, in4091, 
	in4092, in137, in4090, in4089, in4087, in4088, in1694, in1691, 
	in1690, in1689, in372, in369, in292, in289, in562, in245, 
	in552, in556, in559, in386, in132, in23, in80, in25, 
	in81, in79, in82, in24, in26, in86, in88, in87, 
	in83, in34, in4115, in135, in3717, in3724, in141, in2358, 
	in31, in27, in545, in549, in3173, in136, in1, in373, 
	in145, in2824, in140,
	out658, out690, out767, out807, out654, out651, out648, 
	out645, out642, out670, out667, out664, out661, out688, out685, 
	out682, out679, out676, out702, out699, out696, out693, out727, 
	out732, out737, out742, out747, out752, out757, out762, out722, 
	out712, out772, out777, out782, out787, out792, out797, out802, 
	out859, out824, out826, out832, out828, out830, out834, out836, 
	out838, out822, out863, out871, out865, out867, out869, out873, 
	out875, out877, out861, out629, out591, out618, out615, out621, 
	out588, out626, out632, out843, out882, out585, out575, out598, 
	out610, out998, out1002, out1000, out1004, out854, out623, out813, 
	out818, out707, out715, out639, out673, out636, out820, out717, 
	out704, out593, out594, out602, out809, out611, out599, out612, 
	out600, out850, out848, out849, out851, out887, out298, out926, 
	out892, out973, out993, out144, out601, out847, out815, out634, 
	out810, out845, out656, out923, out939, out921, out978, out949, 
	out889, out603, out604, out606);

   input
	in293, in302, in308, in316, in324, in341, in351, 
	in361, in299, in307, in315, in323, in331, in338, in348, 
	in358, in366, in206, in210, in218, in226, in234, in257, 
	in265, in273, in281, in209, in217, in225, in233, in241, 
	in264, in272, in280, in288, in54, in4, in2174, in1497, 
	in332, in335, in479, in490, in503, in514, in523, in534, 
	in446, in457, in468, in422, in435, in389, in400, in411, 
	in374, in191, in200, in194, in197, in203, in149, in155, 
	in188, in182, in161, in170, in164, in167, in173, in146, 
	in152, in158, in185, in109, in43, in46, in100, in91, 
	in76, in73, in67, in11, in106, in37, in49, in103, 
	in40, in20, in17, in70, in61, in123, in52, in121, 
	in116, in112, in130, in119, in129, in131, in115, in122, 
	in114, in53, in113, in128, in127, in126, in117, in176, 
	in179, in14, in64, in248, in251, in242, in254, in3552, 
	in3550, in3546, in3548, in120, in94, in118, in97, in4091, 
	in4092, in137, in4090, in4089, in4087, in4088, in1694, in1691, 
	in1690, in1689, in372, in369, in292, in289, in562, in245, 
	in552, in556, in559, in386, in132, in23, in80, in25, 
	in81, in79, in82, in24, in26, in86, in88, in87, 
	in83, in34, in4115, in135, in3717, in3724, in141, in2358, 
	in31, in27, in545, in549, in3173, in136, in1, in373, 
	in145, in2824, in140;

   output
	out658, out690, out767, out807, out654, out651, out648, 
	out645, out642, out670, out667, out664, out661, out688, out685, 
	out682, out679, out676, out702, out699, out696, out693, out727, 
	out732, out737, out742, out747, out752, out757, out762, out722, 
	out712, out772, out777, out782, out787, out792, out797, out802, 
	out859, out824, out826, out832, out828, out830, out834, out836, 
	out838, out822, out863, out871, out865, out867, out869, out873, 
	out875, out877, out861, out629, out591, out618, out615, out621, 
	out588, out626, out632, out843, out882, out585, out575, out598, 
	out610, out998, out1002, out1000, out1004, out854, out623, out813, 
	out818, out707, out715, out639, out673, out636, out820, out717, 
	out704, out593, out594, out602, out809, out611, out599, out612, 
	out600, out850, out848, out849, out851, out887, out298, out926, 
	out892, out973, out993, out144, out601, out847, out815, out634, 
	out810, out845, out656, out923, out939, out921, out978, out949, 
	out889, out603, out604, out606;

inv M1_Mux9_0_Mux4_0_Mux2_0(in332, M1_Mux9_0_Mux4_0_Not_ContIn);
and2 M1_Mux9_0_Mux4_0_Mux2_1(in361, M1_Mux9_0_Mux4_0_Not_ContIn, M1_Mux9_0_Mux4_0_line1);
and2 M1_Mux9_0_Mux4_0_Mux2_2(in366, in332, M1_Mux9_0_Mux4_0_line2);
or2 M1_Mux9_0_Mux4_0_Mux2_3(M1_Mux9_0_Mux4_0_line1, M1_Mux9_0_Mux4_0_line2, Xbus_0);
inv M1_Mux9_0_Mux4_1_Mux2_0(in332, M1_Mux9_0_Mux4_1_Not_ContIn);
and2 M1_Mux9_0_Mux4_1_Mux2_1(in351, M1_Mux9_0_Mux4_1_Not_ContIn, M1_Mux9_0_Mux4_1_line1);
and2 M1_Mux9_0_Mux4_1_Mux2_2(in358, in332, M1_Mux9_0_Mux4_1_line2);
or2 M1_Mux9_0_Mux4_1_Mux2_3(M1_Mux9_0_Mux4_1_line1, M1_Mux9_0_Mux4_1_line2, Xbus_1);
inv M1_Mux9_0_Mux4_2_Mux2_0(in332, M1_Mux9_0_Mux4_2_Not_ContIn);
and2 M1_Mux9_0_Mux4_2_Mux2_1(in341, M1_Mux9_0_Mux4_2_Not_ContIn, M1_Mux9_0_Mux4_2_line1);
and2 M1_Mux9_0_Mux4_2_Mux2_2(in348, in332, M1_Mux9_0_Mux4_2_line2);
or2 M1_Mux9_0_Mux4_2_Mux2_3(M1_Mux9_0_Mux4_2_line1, M1_Mux9_0_Mux4_2_line2, Xbus_2);
inv M1_Mux9_0_Mux4_3_Mux2_0(in332, M1_Mux9_0_Mux4_3_Not_ContIn);
and2 M1_Mux9_0_Mux4_3_Mux2_1(vdd, M1_Mux9_0_Mux4_3_Not_ContIn, M1_Mux9_0_Mux4_3_line1);
and2 M1_Mux9_0_Mux4_3_Mux2_2(in338, in332, M1_Mux9_0_Mux4_3_line2);
or2 M1_Mux9_0_Mux4_3_Mux2_3(M1_Mux9_0_Mux4_3_line1, M1_Mux9_0_Mux4_3_line2, Xbus_3);
inv M1_Mux9_1_Mux4_0_Mux2_0(in332, M1_Mux9_1_Mux4_0_Not_ContIn);
and2 M1_Mux9_1_Mux4_0_Mux2_1(in324, M1_Mux9_1_Mux4_0_Not_ContIn, M1_Mux9_1_Mux4_0_line1);
and2 M1_Mux9_1_Mux4_0_Mux2_2(in331, in332, M1_Mux9_1_Mux4_0_line2);
or2 M1_Mux9_1_Mux4_0_Mux2_3(M1_Mux9_1_Mux4_0_line1, M1_Mux9_1_Mux4_0_line2, Xbus_4);
inv M1_Mux9_1_Mux4_1_Mux2_0(in332, M1_Mux9_1_Mux4_1_Not_ContIn);
and2 M1_Mux9_1_Mux4_1_Mux2_1(in316, M1_Mux9_1_Mux4_1_Not_ContIn, M1_Mux9_1_Mux4_1_line1);
and2 M1_Mux9_1_Mux4_1_Mux2_2(in323, in332, M1_Mux9_1_Mux4_1_line2);
or2 M1_Mux9_1_Mux4_1_Mux2_3(M1_Mux9_1_Mux4_1_line1, M1_Mux9_1_Mux4_1_line2, Xbus_5);
inv M1_Mux9_1_Mux4_2_Mux2_0(in332, M1_Mux9_1_Mux4_2_Not_ContIn);
and2 M1_Mux9_1_Mux4_2_Mux2_1(in308, M1_Mux9_1_Mux4_2_Not_ContIn, M1_Mux9_1_Mux4_2_line1);
and2 M1_Mux9_1_Mux4_2_Mux2_2(in315, in332, M1_Mux9_1_Mux4_2_line2);
or2 M1_Mux9_1_Mux4_2_Mux2_3(M1_Mux9_1_Mux4_2_line1, M1_Mux9_1_Mux4_2_line2, Xbus_6);
inv M1_Mux9_1_Mux4_3_Mux2_0(in332, M1_Mux9_1_Mux4_3_Not_ContIn);
and2 M1_Mux9_1_Mux4_3_Mux2_1(in302, M1_Mux9_1_Mux4_3_Not_ContIn, M1_Mux9_1_Mux4_3_line1);
and2 M1_Mux9_1_Mux4_3_Mux2_2(in307, in332, M1_Mux9_1_Mux4_3_line2);
or2 M1_Mux9_1_Mux4_3_Mux2_3(M1_Mux9_1_Mux4_3_line1, M1_Mux9_1_Mux4_3_line2, Xbus_7);
inv M1_Mux9_2_Mux2_0(in332, M1_Mux9_2_Not_ContIn);
and2 M1_Mux9_2_Mux2_1(in293, M1_Mux9_2_Not_ContIn, M1_Mux9_2_line1);
and2 M1_Mux9_2_Mux2_2(in299, in332, M1_Mux9_2_line2);
or2 M1_Mux9_2_Mux2_3(M1_Mux9_2_line1, M1_Mux9_2_line2, Xbus_8);
inv M2_Mux9_0_Mux4_0_Mux2_0(in335, M2_Mux9_0_Mux4_0_Not_ContIn);
and2 M2_Mux9_0_Mux4_0_Mux2_1(in281, M2_Mux9_0_Mux4_0_Not_ContIn, M2_Mux9_0_Mux4_0_line1);
and2 M2_Mux9_0_Mux4_0_Mux2_2(in288, in335, M2_Mux9_0_Mux4_0_line2);
or2 M2_Mux9_0_Mux4_0_Mux2_3(M2_Mux9_0_Mux4_0_line1, M2_Mux9_0_Mux4_0_line2, Ybus_0);
inv M2_Mux9_0_Mux4_1_Mux2_0(in335, M2_Mux9_0_Mux4_1_Not_ContIn);
and2 M2_Mux9_0_Mux4_1_Mux2_1(in273, M2_Mux9_0_Mux4_1_Not_ContIn, M2_Mux9_0_Mux4_1_line1);
and2 M2_Mux9_0_Mux4_1_Mux2_2(in280, in335, M2_Mux9_0_Mux4_1_line2);
or2 M2_Mux9_0_Mux4_1_Mux2_3(M2_Mux9_0_Mux4_1_line1, M2_Mux9_0_Mux4_1_line2, Ybus_1);
inv M2_Mux9_0_Mux4_2_Mux2_0(in335, M2_Mux9_0_Mux4_2_Not_ContIn);
and2 M2_Mux9_0_Mux4_2_Mux2_1(in265, M2_Mux9_0_Mux4_2_Not_ContIn, M2_Mux9_0_Mux4_2_line1);
and2 M2_Mux9_0_Mux4_2_Mux2_2(in272, in335, M2_Mux9_0_Mux4_2_line2);
or2 M2_Mux9_0_Mux4_2_Mux2_3(M2_Mux9_0_Mux4_2_line1, M2_Mux9_0_Mux4_2_line2, Ybus_2);
inv M2_Mux9_0_Mux4_3_Mux2_0(in335, M2_Mux9_0_Mux4_3_Not_ContIn);
and2 M2_Mux9_0_Mux4_3_Mux2_1(in257, M2_Mux9_0_Mux4_3_Not_ContIn, M2_Mux9_0_Mux4_3_line1);
and2 M2_Mux9_0_Mux4_3_Mux2_2(in264, in335, M2_Mux9_0_Mux4_3_line2);
or2 M2_Mux9_0_Mux4_3_Mux2_3(M2_Mux9_0_Mux4_3_line1, M2_Mux9_0_Mux4_3_line2, Ybus_3);
inv M2_Mux9_1_Mux4_0_Mux2_0(in335, M2_Mux9_1_Mux4_0_Not_ContIn);
and2 M2_Mux9_1_Mux4_0_Mux2_1(in234, M2_Mux9_1_Mux4_0_Not_ContIn, M2_Mux9_1_Mux4_0_line1);
and2 M2_Mux9_1_Mux4_0_Mux2_2(in241, in335, M2_Mux9_1_Mux4_0_line2);
or2 M2_Mux9_1_Mux4_0_Mux2_3(M2_Mux9_1_Mux4_0_line1, M2_Mux9_1_Mux4_0_line2, Ybus_4);
inv M2_Mux9_1_Mux4_1_Mux2_0(in335, M2_Mux9_1_Mux4_1_Not_ContIn);
and2 M2_Mux9_1_Mux4_1_Mux2_1(in226, M2_Mux9_1_Mux4_1_Not_ContIn, M2_Mux9_1_Mux4_1_line1);
and2 M2_Mux9_1_Mux4_1_Mux2_2(in233, in335, M2_Mux9_1_Mux4_1_line2);
or2 M2_Mux9_1_Mux4_1_Mux2_3(M2_Mux9_1_Mux4_1_line1, M2_Mux9_1_Mux4_1_line2, Ybus_5);
inv M2_Mux9_1_Mux4_2_Mux2_0(in335, M2_Mux9_1_Mux4_2_Not_ContIn);
and2 M2_Mux9_1_Mux4_2_Mux2_1(in218, M2_Mux9_1_Mux4_2_Not_ContIn, M2_Mux9_1_Mux4_2_line1);
and2 M2_Mux9_1_Mux4_2_Mux2_2(in225, in335, M2_Mux9_1_Mux4_2_line2);
or2 M2_Mux9_1_Mux4_2_Mux2_3(M2_Mux9_1_Mux4_2_line1, M2_Mux9_1_Mux4_2_line2, Ybus_6);
inv M2_Mux9_1_Mux4_3_Mux2_0(in335, M2_Mux9_1_Mux4_3_Not_ContIn);
and2 M2_Mux9_1_Mux4_3_Mux2_1(in210, M2_Mux9_1_Mux4_3_Not_ContIn, M2_Mux9_1_Mux4_3_line1);
and2 M2_Mux9_1_Mux4_3_Mux2_2(in217, in335, M2_Mux9_1_Mux4_3_line2);
or2 M2_Mux9_1_Mux4_3_Mux2_3(M2_Mux9_1_Mux4_3_line1, M2_Mux9_1_Mux4_3_line2, Ybus_7);
inv M2_Mux9_2_Mux2_0(in335, M2_Mux9_2_Not_ContIn);
and2 M2_Mux9_2_Mux2_1(in206, M2_Mux9_2_Not_ContIn, M2_Mux9_2_line1);
and2 M2_Mux9_2_Mux2_2(in209, in335, M2_Mux9_2_line2);
or2 M2_Mux9_2_Mux2_3(M2_Mux9_2_line1, M2_Mux9_2_line2, Ybus_8);
inv M3_CalP0_LP0_CL0_LB0_Mux2_0(in361, M3_CalP0_LP0_CL0_LB0_Not_ContIn);
and2 M3_CalP0_LP0_CL0_LB0_Mux2_1(in254, M3_CalP0_LP0_CL0_LB0_Not_ContIn, M3_CalP0_LP0_CL0_LB0_line1);
and2 M3_CalP0_LP0_CL0_LB0_Mux2_2(in242, in361, M3_CalP0_LP0_CL0_LB0_line2);
or2 M3_CalP0_LP0_CL0_LB0_Mux2_3(M3_CalP0_LP0_CL0_LB0_line1, M3_CalP0_LP0_CL0_LB0_line2, M3_CalP0_LP0_CL0_line0);
inv M3_CalP0_LP0_CL0_LB1_Mux2_0(in361, M3_CalP0_LP0_CL0_LB1_Not_ContIn);
and2 M3_CalP0_LP0_CL0_LB1_Mux2_1(in251, M3_CalP0_LP0_CL0_LB1_Not_ContIn, M3_CalP0_LP0_CL0_LB1_line1);
and2 M3_CalP0_LP0_CL0_LB1_Mux2_2(in248, in361, M3_CalP0_LP0_CL0_LB1_line2);
or2 M3_CalP0_LP0_CL0_LB1_Mux2_3(M3_CalP0_LP0_CL0_LB1_line1, M3_CalP0_LP0_CL0_LB1_line2, M3_CalP0_LP0_CL0_line1);
or2 M3_CalP0_LP0_CL0_LB2(vdd, M3_CalP0_LP0_CL0_line0, M3_CalP0_LP0_CL0_line2);
nand2 M3_CalP0_LP0_CL0_LB3(vdd, M3_CalP0_LP0_CL0_line1, M3_CalP0_LP0_CL0_line3);
and2 M3_CalP0_LP0_CL0_LB4(M3_CalP0_LP0_CL0_line2, M3_CalP0_LP0_CL0_line3, M3_CalP0_LogicOut_0);
inv M3_CalP0_LP0_CL1_LB0_Mux2_0(in351, M3_CalP0_LP0_CL1_LB0_Not_ContIn);
and2 M3_CalP0_LP0_CL1_LB0_Mux2_1(in254, M3_CalP0_LP0_CL1_LB0_Not_ContIn, M3_CalP0_LP0_CL1_LB0_line1);
and2 M3_CalP0_LP0_CL1_LB0_Mux2_2(in242, in351, M3_CalP0_LP0_CL1_LB0_line2);
or2 M3_CalP0_LP0_CL1_LB0_Mux2_3(M3_CalP0_LP0_CL1_LB0_line1, M3_CalP0_LP0_CL1_LB0_line2, M3_CalP0_LP0_CL1_line0);
inv M3_CalP0_LP0_CL1_LB1_Mux2_0(in351, M3_CalP0_LP0_CL1_LB1_Not_ContIn);
and2 M3_CalP0_LP0_CL1_LB1_Mux2_1(in251, M3_CalP0_LP0_CL1_LB1_Not_ContIn, M3_CalP0_LP0_CL1_LB1_line1);
and2 M3_CalP0_LP0_CL1_LB1_Mux2_2(in248, in351, M3_CalP0_LP0_CL1_LB1_line2);
or2 M3_CalP0_LP0_CL1_LB1_Mux2_3(M3_CalP0_LP0_CL1_LB1_line1, M3_CalP0_LP0_CL1_LB1_line2, M3_CalP0_LP0_CL1_line1);
or2 M3_CalP0_LP0_CL1_LB2(in534, M3_CalP0_LP0_CL1_line0, M3_CalP0_LP0_CL1_line2);
nand2 M3_CalP0_LP0_CL1_LB3(in534, M3_CalP0_LP0_CL1_line1, M3_CalP0_LP0_CL1_line3);
and2 M3_CalP0_LP0_CL1_LB4(M3_CalP0_LP0_CL1_line2, M3_CalP0_LP0_CL1_line3, M3_CalP0_LogicOut_1);
inv M3_CalP0_LP0_CL2_LB0_Mux2_0(in341, M3_CalP0_LP0_CL2_LB0_Not_ContIn);
and2 M3_CalP0_LP0_CL2_LB0_Mux2_1(in254, M3_CalP0_LP0_CL2_LB0_Not_ContIn, M3_CalP0_LP0_CL2_LB0_line1);
and2 M3_CalP0_LP0_CL2_LB0_Mux2_2(in242, in341, M3_CalP0_LP0_CL2_LB0_line2);
or2 M3_CalP0_LP0_CL2_LB0_Mux2_3(M3_CalP0_LP0_CL2_LB0_line1, M3_CalP0_LP0_CL2_LB0_line2, M3_CalP0_LP0_CL2_line0);
inv M3_CalP0_LP0_CL2_LB1_Mux2_0(in341, M3_CalP0_LP0_CL2_LB1_Not_ContIn);
and2 M3_CalP0_LP0_CL2_LB1_Mux2_1(in251, M3_CalP0_LP0_CL2_LB1_Not_ContIn, M3_CalP0_LP0_CL2_LB1_line1);
and2 M3_CalP0_LP0_CL2_LB1_Mux2_2(in248, in341, M3_CalP0_LP0_CL2_LB1_line2);
or2 M3_CalP0_LP0_CL2_LB1_Mux2_3(M3_CalP0_LP0_CL2_LB1_line1, M3_CalP0_LP0_CL2_LB1_line2, M3_CalP0_LP0_CL2_line1);
or2 M3_CalP0_LP0_CL2_LB2(in523, M3_CalP0_LP0_CL2_line0, M3_CalP0_LP0_CL2_line2);
nand2 M3_CalP0_LP0_CL2_LB3(in523, M3_CalP0_LP0_CL2_line1, M3_CalP0_LP0_CL2_line3);
and2 M3_CalP0_LP0_CL2_LB4(M3_CalP0_LP0_CL2_line2, M3_CalP0_LP0_CL2_line3, M3_CalP0_LogicOut_2);
inv M3_CalP0_LP0_CL3_LB0_Mux2_0(vdd, M3_CalP0_LP0_CL3_LB0_Not_ContIn);
and2 M3_CalP0_LP0_CL3_LB0_Mux2_1(in254, M3_CalP0_LP0_CL3_LB0_Not_ContIn, M3_CalP0_LP0_CL3_LB0_line1);
and2 M3_CalP0_LP0_CL3_LB0_Mux2_2(in242, vdd, M3_CalP0_LP0_CL3_LB0_line2);
or2 M3_CalP0_LP0_CL3_LB0_Mux2_3(M3_CalP0_LP0_CL3_LB0_line1, M3_CalP0_LP0_CL3_LB0_line2, M3_CalP0_LP0_CL3_line0);
inv M3_CalP0_LP0_CL3_LB1_Mux2_0(vdd, M3_CalP0_LP0_CL3_LB1_Not_ContIn);
and2 M3_CalP0_LP0_CL3_LB1_Mux2_1(in251, M3_CalP0_LP0_CL3_LB1_Not_ContIn, M3_CalP0_LP0_CL3_LB1_line1);
and2 M3_CalP0_LP0_CL3_LB1_Mux2_2(in248, vdd, M3_CalP0_LP0_CL3_LB1_line2);
or2 M3_CalP0_LP0_CL3_LB1_Mux2_3(M3_CalP0_LP0_CL3_LB1_line1, M3_CalP0_LP0_CL3_LB1_line2, M3_CalP0_LP0_CL3_line1);
or2 M3_CalP0_LP0_CL3_LB2(in514, M3_CalP0_LP0_CL3_line0, M3_CalP0_LP0_CL3_line2);
nand2 M3_CalP0_LP0_CL3_LB3(in514, M3_CalP0_LP0_CL3_line1, M3_CalP0_LP0_CL3_line3);
and2 M3_CalP0_LP0_CL3_LB4(M3_CalP0_LP0_CL3_line2, M3_CalP0_LP0_CL3_line3, M3_CalP0_LogicOut_3);
inv M3_CalP0_LP0_CL4_LB0_Mux2_0(in324, M3_CalP0_LP0_CL4_LB0_Not_ContIn);
and2 M3_CalP0_LP0_CL4_LB0_Mux2_1(in254, M3_CalP0_LP0_CL4_LB0_Not_ContIn, M3_CalP0_LP0_CL4_LB0_line1);
and2 M3_CalP0_LP0_CL4_LB0_Mux2_2(in242, in324, M3_CalP0_LP0_CL4_LB0_line2);
or2 M3_CalP0_LP0_CL4_LB0_Mux2_3(M3_CalP0_LP0_CL4_LB0_line1, M3_CalP0_LP0_CL4_LB0_line2, M3_CalP0_LP0_CL4_line0);
inv M3_CalP0_LP0_CL4_LB1_Mux2_0(in324, M3_CalP0_LP0_CL4_LB1_Not_ContIn);
and2 M3_CalP0_LP0_CL4_LB1_Mux2_1(in251, M3_CalP0_LP0_CL4_LB1_Not_ContIn, M3_CalP0_LP0_CL4_LB1_line1);
and2 M3_CalP0_LP0_CL4_LB1_Mux2_2(in248, in324, M3_CalP0_LP0_CL4_LB1_line2);
or2 M3_CalP0_LP0_CL4_LB1_Mux2_3(M3_CalP0_LP0_CL4_LB1_line1, M3_CalP0_LP0_CL4_LB1_line2, M3_CalP0_LP0_CL4_line1);
or2 M3_CalP0_LP0_CL4_LB2(in503, M3_CalP0_LP0_CL4_line0, M3_CalP0_LP0_CL4_line2);
nand2 M3_CalP0_LP0_CL4_LB3(in503, M3_CalP0_LP0_CL4_line1, M3_CalP0_LP0_CL4_line3);
and2 M3_CalP0_LP0_CL4_LB4(M3_CalP0_LP0_CL4_line2, M3_CalP0_LP0_CL4_line3, M3_CalP0_LogicOut_4);
inv M3_CalP0_LP0_CL5_LB0_Mux2_0(in316, M3_CalP0_LP0_CL5_LB0_Not_ContIn);
and2 M3_CalP0_LP0_CL5_LB0_Mux2_1(in254, M3_CalP0_LP0_CL5_LB0_Not_ContIn, M3_CalP0_LP0_CL5_LB0_line1);
and2 M3_CalP0_LP0_CL5_LB0_Mux2_2(in242, in316, M3_CalP0_LP0_CL5_LB0_line2);
or2 M3_CalP0_LP0_CL5_LB0_Mux2_3(M3_CalP0_LP0_CL5_LB0_line1, M3_CalP0_LP0_CL5_LB0_line2, M3_CalP0_LP0_CL5_line0);
inv M3_CalP0_LP0_CL5_LB1_Mux2_0(in316, M3_CalP0_LP0_CL5_LB1_Not_ContIn);
and2 M3_CalP0_LP0_CL5_LB1_Mux2_1(in251, M3_CalP0_LP0_CL5_LB1_Not_ContIn, M3_CalP0_LP0_CL5_LB1_line1);
and2 M3_CalP0_LP0_CL5_LB1_Mux2_2(in248, in316, M3_CalP0_LP0_CL5_LB1_line2);
or2 M3_CalP0_LP0_CL5_LB1_Mux2_3(M3_CalP0_LP0_CL5_LB1_line1, M3_CalP0_LP0_CL5_LB1_line2, M3_CalP0_LP0_CL5_line1);
or2 M3_CalP0_LP0_CL5_LB2(in490, M3_CalP0_LP0_CL5_line0, M3_CalP0_LP0_CL5_line2);
nand2 M3_CalP0_LP0_CL5_LB3(in490, M3_CalP0_LP0_CL5_line1, M3_CalP0_LP0_CL5_line3);
and2 M3_CalP0_LP0_CL5_LB4(M3_CalP0_LP0_CL5_line2, M3_CalP0_LP0_CL5_line3, M3_CalP0_LogicOut_5);
inv M3_CalP0_LP0_CL6_LB0_Mux2_0(in308, M3_CalP0_LP0_CL6_LB0_Not_ContIn);
and2 M3_CalP0_LP0_CL6_LB0_Mux2_1(in254, M3_CalP0_LP0_CL6_LB0_Not_ContIn, M3_CalP0_LP0_CL6_LB0_line1);
and2 M3_CalP0_LP0_CL6_LB0_Mux2_2(in242, in308, M3_CalP0_LP0_CL6_LB0_line2);
or2 M3_CalP0_LP0_CL6_LB0_Mux2_3(M3_CalP0_LP0_CL6_LB0_line1, M3_CalP0_LP0_CL6_LB0_line2, M3_CalP0_LP0_CL6_line0);
inv M3_CalP0_LP0_CL6_LB1_Mux2_0(in308, M3_CalP0_LP0_CL6_LB1_Not_ContIn);
and2 M3_CalP0_LP0_CL6_LB1_Mux2_1(in251, M3_CalP0_LP0_CL6_LB1_Not_ContIn, M3_CalP0_LP0_CL6_LB1_line1);
and2 M3_CalP0_LP0_CL6_LB1_Mux2_2(in248, in308, M3_CalP0_LP0_CL6_LB1_line2);
or2 M3_CalP0_LP0_CL6_LB1_Mux2_3(M3_CalP0_LP0_CL6_LB1_line1, M3_CalP0_LP0_CL6_LB1_line2, M3_CalP0_LP0_CL6_line1);
or2 M3_CalP0_LP0_CL6_LB2(in479, M3_CalP0_LP0_CL6_line0, M3_CalP0_LP0_CL6_line2);
nand2 M3_CalP0_LP0_CL6_LB3(in479, M3_CalP0_LP0_CL6_line1, M3_CalP0_LP0_CL6_line3);
and2 M3_CalP0_LP0_CL6_LB4(M3_CalP0_LP0_CL6_line2, M3_CalP0_LP0_CL6_line3, M3_CalP0_LogicOut_6);
inv M3_CalP0_LP0_CL7_LB0_Mux2_0(in302, M3_CalP0_LP0_CL7_LB0_Not_ContIn);
and2 M3_CalP0_LP0_CL7_LB0_Mux2_1(in254, M3_CalP0_LP0_CL7_LB0_Not_ContIn, M3_CalP0_LP0_CL7_LB0_line1);
and2 M3_CalP0_LP0_CL7_LB0_Mux2_2(in242, in302, M3_CalP0_LP0_CL7_LB0_line2);
or2 M3_CalP0_LP0_CL7_LB0_Mux2_3(M3_CalP0_LP0_CL7_LB0_line1, M3_CalP0_LP0_CL7_LB0_line2, M3_CalP0_LP0_CL7_line0);
inv M3_CalP0_LP0_CL7_LB1_Mux2_0(in302, M3_CalP0_LP0_CL7_LB1_Not_ContIn);
and2 M3_CalP0_LP0_CL7_LB1_Mux2_1(in251, M3_CalP0_LP0_CL7_LB1_Not_ContIn, M3_CalP0_LP0_CL7_LB1_line1);
and2 M3_CalP0_LP0_CL7_LB1_Mux2_2(in248, in302, M3_CalP0_LP0_CL7_LB1_line2);
or2 M3_CalP0_LP0_CL7_LB1_Mux2_3(M3_CalP0_LP0_CL7_LB1_line1, M3_CalP0_LP0_CL7_LB1_line2, M3_CalP0_LP0_CL7_line1);
or2 M3_CalP0_LP0_CL7_LB2(vdd, M3_CalP0_LP0_CL7_line0, M3_CalP0_LP0_CL7_line2);
nand2 M3_CalP0_LP0_CL7_LB3(vdd, M3_CalP0_LP0_CL7_line1, M3_CalP0_LP0_CL7_line3);
and2 M3_CalP0_LP0_CL7_LB4(M3_CalP0_LP0_CL7_line2, M3_CalP0_LP0_CL7_line3, M3_CalP0_LogicOut_7);
inv M3_CalP0_LP0_CL8_LB0_Mux2_0(in293, M3_CalP0_LP0_CL8_LB0_Not_ContIn);
and2 M3_CalP0_LP0_CL8_LB0_Mux2_1(in254, M3_CalP0_LP0_CL8_LB0_Not_ContIn, M3_CalP0_LP0_CL8_LB0_line1);
and2 M3_CalP0_LP0_CL8_LB0_Mux2_2(in242, in293, M3_CalP0_LP0_CL8_LB0_line2);
or2 M3_CalP0_LP0_CL8_LB0_Mux2_3(M3_CalP0_LP0_CL8_LB0_line1, M3_CalP0_LP0_CL8_LB0_line2, M3_CalP0_LP0_CL8_line0);
inv M3_CalP0_LP0_CL8_LB1_Mux2_0(in293, M3_CalP0_LP0_CL8_LB1_Not_ContIn);
and2 M3_CalP0_LP0_CL8_LB1_Mux2_1(in251, M3_CalP0_LP0_CL8_LB1_Not_ContIn, M3_CalP0_LP0_CL8_LB1_line1);
and2 M3_CalP0_LP0_CL8_LB1_Mux2_2(in248, in293, M3_CalP0_LP0_CL8_LB1_line2);
or2 M3_CalP0_LP0_CL8_LB1_Mux2_3(M3_CalP0_LP0_CL8_LB1_line1, M3_CalP0_LP0_CL8_LB1_line2, M3_CalP0_LP0_CL8_line1);
or2 M3_CalP0_LP0_CL8_LB2(gnd, M3_CalP0_LP0_CL8_line0, M3_CalP0_LP0_CL8_line2);
nand2 M3_CalP0_LP0_CL8_LB3(gnd, M3_CalP0_LP0_CL8_line1, M3_CalP0_LP0_CL8_line3);
and2 M3_CalP0_LP0_CL8_LB4(M3_CalP0_LP0_CL8_line2, M3_CalP0_LP0_CL8_line3, M3_CalP0_LogicOut_8);
inv M3_CalP0_LP1_PT1_Xo0(M3_CalP0_LogicOut_5, M3_CalP0_LP1_PT1_NotA);
inv M3_CalP0_LP1_PT1_Xo1(M3_CalP0_LogicOut_6, M3_CalP0_LP1_PT1_NotB);
nand2 M3_CalP0_LP1_PT1_Xo2(M3_CalP0_LP1_PT1_NotA, M3_CalP0_LogicOut_6, M3_CalP0_LP1_PT1_line2);
nand2 M3_CalP0_LP1_PT1_Xo3(M3_CalP0_LP1_PT1_NotB, M3_CalP0_LogicOut_5, M3_CalP0_LP1_PT1_line3);
nand2 M3_CalP0_LP1_PT1_Xo4(M3_CalP0_LP1_PT1_line2, M3_CalP0_LP1_PT1_line3, M3_CalP0_LP1_line1);
inv M3_CalP0_LP1_PT2_Xo0(M3_CalP0_LogicOut_7, M3_CalP0_LP1_PT2_NotA);
inv M3_CalP0_LP1_PT2_Xo1(M3_CalP0_LogicOut_8, M3_CalP0_LP1_PT2_NotB);
nand2 M3_CalP0_LP1_PT2_Xo2(M3_CalP0_LP1_PT2_NotA, M3_CalP0_LogicOut_8, M3_CalP0_LP1_PT2_line2);
nand2 M3_CalP0_LP1_PT2_Xo3(M3_CalP0_LP1_PT2_NotB, M3_CalP0_LogicOut_7, M3_CalP0_LP1_PT2_line3);
nand2 M3_CalP0_LP1_PT2_Xo4(M3_CalP0_LP1_PT2_line2, M3_CalP0_LP1_PT2_line3, M3_CalP0_LP1_line2);
inv M3_CalP0_LP1_PT3_Xo0(M3_CalP0_LogicOut_1, M3_CalP0_LP1_PT3_NotA);
inv M3_CalP0_LP1_PT3_Xo1(M3_CalP0_LogicOut_2, M3_CalP0_LP1_PT3_NotB);
nand2 M3_CalP0_LP1_PT3_Xo2(M3_CalP0_LP1_PT3_NotA, M3_CalP0_LogicOut_2, M3_CalP0_LP1_PT3_line2);
nand2 M3_CalP0_LP1_PT3_Xo3(M3_CalP0_LP1_PT3_NotB, M3_CalP0_LogicOut_1, M3_CalP0_LP1_PT3_line3);
nand2 M3_CalP0_LP1_PT3_Xo4(M3_CalP0_LP1_PT3_line2, M3_CalP0_LP1_PT3_line3, M3_CalP0_LP1_line3);
inv M3_CalP0_LP1_PT4_Xo0(M3_CalP0_LogicOut_3, M3_CalP0_LP1_PT4_NotA);
inv M3_CalP0_LP1_PT4_Xo1(M3_CalP0_LogicOut_4, M3_CalP0_LP1_PT4_NotB);
nand2 M3_CalP0_LP1_PT4_Xo2(M3_CalP0_LP1_PT4_NotA, M3_CalP0_LogicOut_4, M3_CalP0_LP1_PT4_line2);
nand2 M3_CalP0_LP1_PT4_Xo3(M3_CalP0_LP1_PT4_NotB, M3_CalP0_LogicOut_3, M3_CalP0_LP1_PT4_line3);
nand2 M3_CalP0_LP1_PT4_Xo4(M3_CalP0_LP1_PT4_line2, M3_CalP0_LP1_PT4_line3, M3_CalP0_LP1_line4);
inv M3_CalP0_LP1_PT5_Xo0(M3_CalP0_LP1_line1, M3_CalP0_LP1_PT5_NotA);
inv M3_CalP0_LP1_PT5_Xo1(M3_CalP0_LP1_line2, M3_CalP0_LP1_PT5_NotB);
nand2 M3_CalP0_LP1_PT5_Xo2(M3_CalP0_LP1_PT5_NotA, M3_CalP0_LP1_line2, M3_CalP0_LP1_PT5_line2);
nand2 M3_CalP0_LP1_PT5_Xo3(M3_CalP0_LP1_PT5_NotB, M3_CalP0_LP1_line1, M3_CalP0_LP1_PT5_line3);
nand2 M3_CalP0_LP1_PT5_Xo4(M3_CalP0_LP1_PT5_line2, M3_CalP0_LP1_PT5_line3, M3_CalP0_LP1_line5);
inv M3_CalP0_LP1_PT6_Xo3_0(M3_CalP0_LP1_line3, M3_CalP0_LP1_PT6_NotA);
inv M3_CalP0_LP1_PT6_Xo3_1(M3_CalP0_LogicOut_0, M3_CalP0_LP1_PT6_NotB);
inv M3_CalP0_LP1_PT6_Xo3_2(M3_CalP0_LP1_line4, M3_CalP0_LP1_PT6_NotC);
and3 M3_CalP0_LP1_PT6_Xo3_3(M3_CalP0_LP1_PT6_NotA, M3_CalP0_LP1_PT6_NotB, M3_CalP0_LP1_line4, M3_CalP0_LP1_PT6_line3);
and3 M3_CalP0_LP1_PT6_Xo3_4(M3_CalP0_LP1_PT6_NotA, M3_CalP0_LogicOut_0, M3_CalP0_LP1_PT6_NotC, M3_CalP0_LP1_PT6_line4);
and3 M3_CalP0_LP1_PT6_Xo3_5(M3_CalP0_LP1_line3, M3_CalP0_LP1_PT6_NotB, M3_CalP0_LP1_PT6_NotC, M3_CalP0_LP1_PT6_line5);
and3 M3_CalP0_LP1_PT6_Xo3_6(M3_CalP0_LP1_line3, M3_CalP0_LogicOut_0, M3_CalP0_LP1_line4, M3_CalP0_LP1_PT6_line6);
nor2 M3_CalP0_LP1_PT6_Xo3_7(M3_CalP0_LP1_PT6_line3, M3_CalP0_LP1_PT6_line4, M3_CalP0_LP1_PT6_line7);
nor2 M3_CalP0_LP1_PT6_Xo3_8(M3_CalP0_LP1_PT6_line5, M3_CalP0_LP1_PT6_line6, M3_CalP0_LP1_PT6_line8);
nand2 M3_CalP0_LP1_PT6_Xo3_9(M3_CalP0_LP1_PT6_line7, M3_CalP0_LP1_PT6_line8, M3_CalP0_LP1_line6);
inv M3_CalP0_LP1_PT7_Xo0(M3_CalP0_LP1_line5, M3_CalP0_LP1_PT7_NotA);
inv M3_CalP0_LP1_PT7_Xo1(M3_CalP0_LP1_line6, M3_CalP0_LP1_PT7_NotB);
nand2 M3_CalP0_LP1_PT7_Xo2(M3_CalP0_LP1_PT7_NotA, M3_CalP0_LP1_line6, M3_CalP0_LP1_PT7_line2);
nand2 M3_CalP0_LP1_PT7_Xo3(M3_CalP0_LP1_PT7_NotB, M3_CalP0_LP1_line5, M3_CalP0_LP1_PT7_line3);
nand2 M3_CalP0_LP1_PT7_Xo4(M3_CalP0_LP1_PT7_line2, M3_CalP0_LP1_PT7_line3, M3_LogicPar);
and2 M3_CalP1_SP0_GP9_0(Xbus_0, vdd, M3_CalP1_Genbus_0);
and2 M3_CalP1_SP0_GP9_1(Xbus_1, in534, M3_CalP1_Genbus_1);
and2 M3_CalP1_SP0_GP9_2(Xbus_2, in523, M3_CalP1_Genbus_2);
and2 M3_CalP1_SP0_GP9_3(Xbus_3, in514, M3_CalP1_Genbus_3);
and2 M3_CalP1_SP0_GP9_4(Xbus_4, in503, M3_CalP1_Genbus_4);
and2 M3_CalP1_SP0_GP9_5(Xbus_5, in490, M3_CalP1_Genbus_5);
and2 M3_CalP1_SP0_GP9_6(Xbus_6, in479, M3_CalP1_Genbus_6);
and2 M3_CalP1_SP0_GP9_7(Xbus_7, vdd, M3_CalP1_Genbus_7);
and2 M3_CalP1_SP0_GP9_8(Xbus_8, vdd, M3_CalP1_Genbus_8);
inv M3_CalP1_SP0_GP9_9_Xo0(Xbus_0, M3_CalP1_SP0_GP9_9_NotA);
inv M3_CalP1_SP0_GP9_9_Xo1(vdd, M3_CalP1_SP0_GP9_9_NotB);
nand2 M3_CalP1_SP0_GP9_9_Xo2(M3_CalP1_SP0_GP9_9_NotA, vdd, M3_CalP1_SP0_GP9_9_line2);
nand2 M3_CalP1_SP0_GP9_9_Xo3(M3_CalP1_SP0_GP9_9_NotB, Xbus_0, M3_CalP1_SP0_GP9_9_line3);
nand2 M3_CalP1_SP0_GP9_9_Xo4(M3_CalP1_SP0_GP9_9_line2, M3_CalP1_SP0_GP9_9_line3, M3_CalP1_Propbus_0);
inv M3_CalP1_SP0_GP9_10_Xo0(Xbus_1, M3_CalP1_SP0_GP9_10_NotA);
inv M3_CalP1_SP0_GP9_10_Xo1(in534, M3_CalP1_SP0_GP9_10_NotB);
nand2 M3_CalP1_SP0_GP9_10_Xo2(M3_CalP1_SP0_GP9_10_NotA, in534, M3_CalP1_SP0_GP9_10_line2);
nand2 M3_CalP1_SP0_GP9_10_Xo3(M3_CalP1_SP0_GP9_10_NotB, Xbus_1, M3_CalP1_SP0_GP9_10_line3);
nand2 M3_CalP1_SP0_GP9_10_Xo4(M3_CalP1_SP0_GP9_10_line2, M3_CalP1_SP0_GP9_10_line3, M3_CalP1_Propbus_1);
inv M3_CalP1_SP0_GP9_11_Xo0(Xbus_2, M3_CalP1_SP0_GP9_11_NotA);
inv M3_CalP1_SP0_GP9_11_Xo1(in523, M3_CalP1_SP0_GP9_11_NotB);
nand2 M3_CalP1_SP0_GP9_11_Xo2(M3_CalP1_SP0_GP9_11_NotA, in523, M3_CalP1_SP0_GP9_11_line2);
nand2 M3_CalP1_SP0_GP9_11_Xo3(M3_CalP1_SP0_GP9_11_NotB, Xbus_2, M3_CalP1_SP0_GP9_11_line3);
nand2 M3_CalP1_SP0_GP9_11_Xo4(M3_CalP1_SP0_GP9_11_line2, M3_CalP1_SP0_GP9_11_line3, M3_CalP1_Propbus_2);
inv M3_CalP1_SP0_GP9_12_Xo0(Xbus_3, M3_CalP1_SP0_GP9_12_NotA);
inv M3_CalP1_SP0_GP9_12_Xo1(in514, M3_CalP1_SP0_GP9_12_NotB);
nand2 M3_CalP1_SP0_GP9_12_Xo2(M3_CalP1_SP0_GP9_12_NotA, in514, M3_CalP1_SP0_GP9_12_line2);
nand2 M3_CalP1_SP0_GP9_12_Xo3(M3_CalP1_SP0_GP9_12_NotB, Xbus_3, M3_CalP1_SP0_GP9_12_line3);
nand2 M3_CalP1_SP0_GP9_12_Xo4(M3_CalP1_SP0_GP9_12_line2, M3_CalP1_SP0_GP9_12_line3, M3_CalP1_Propbus_3);
inv M3_CalP1_SP0_GP9_13_Xo0(Xbus_4, M3_CalP1_SP0_GP9_13_NotA);
inv M3_CalP1_SP0_GP9_13_Xo1(in503, M3_CalP1_SP0_GP9_13_NotB);
nand2 M3_CalP1_SP0_GP9_13_Xo2(M3_CalP1_SP0_GP9_13_NotA, in503, M3_CalP1_SP0_GP9_13_line2);
nand2 M3_CalP1_SP0_GP9_13_Xo3(M3_CalP1_SP0_GP9_13_NotB, Xbus_4, M3_CalP1_SP0_GP9_13_line3);
nand2 M3_CalP1_SP0_GP9_13_Xo4(M3_CalP1_SP0_GP9_13_line2, M3_CalP1_SP0_GP9_13_line3, M3_CalP1_Propbus_4);
inv M3_CalP1_SP0_GP9_14_Xo0(Xbus_5, M3_CalP1_SP0_GP9_14_NotA);
inv M3_CalP1_SP0_GP9_14_Xo1(in490, M3_CalP1_SP0_GP9_14_NotB);
nand2 M3_CalP1_SP0_GP9_14_Xo2(M3_CalP1_SP0_GP9_14_NotA, in490, M3_CalP1_SP0_GP9_14_line2);
nand2 M3_CalP1_SP0_GP9_14_Xo3(M3_CalP1_SP0_GP9_14_NotB, Xbus_5, M3_CalP1_SP0_GP9_14_line3);
nand2 M3_CalP1_SP0_GP9_14_Xo4(M3_CalP1_SP0_GP9_14_line2, M3_CalP1_SP0_GP9_14_line3, M3_CalP1_Propbus_5);
inv M3_CalP1_SP0_GP9_15_Xo0(Xbus_6, M3_CalP1_SP0_GP9_15_NotA);
inv M3_CalP1_SP0_GP9_15_Xo1(in479, M3_CalP1_SP0_GP9_15_NotB);
nand2 M3_CalP1_SP0_GP9_15_Xo2(M3_CalP1_SP0_GP9_15_NotA, in479, M3_CalP1_SP0_GP9_15_line2);
nand2 M3_CalP1_SP0_GP9_15_Xo3(M3_CalP1_SP0_GP9_15_NotB, Xbus_6, M3_CalP1_SP0_GP9_15_line3);
nand2 M3_CalP1_SP0_GP9_15_Xo4(M3_CalP1_SP0_GP9_15_line2, M3_CalP1_SP0_GP9_15_line3, M3_CalP1_Propbus_6);
inv M3_CalP1_SP0_GP9_16_Xo0(Xbus_7, M3_CalP1_SP0_GP9_16_NotA);
inv M3_CalP1_SP0_GP9_16_Xo1(vdd, M3_CalP1_SP0_GP9_16_NotB);
nand2 M3_CalP1_SP0_GP9_16_Xo2(M3_CalP1_SP0_GP9_16_NotA, vdd, M3_CalP1_SP0_GP9_16_line2);
nand2 M3_CalP1_SP0_GP9_16_Xo3(M3_CalP1_SP0_GP9_16_NotB, Xbus_7, M3_CalP1_SP0_GP9_16_line3);
nand2 M3_CalP1_SP0_GP9_16_Xo4(M3_CalP1_SP0_GP9_16_line2, M3_CalP1_SP0_GP9_16_line3, M3_CalP1_Propbus_7);
inv M3_CalP1_SP0_GP9_17_Xo0(Xbus_8, M3_CalP1_SP0_GP9_17_NotA);
inv M3_CalP1_SP0_GP9_17_Xo1(vdd, M3_CalP1_SP0_GP9_17_NotB);
nand2 M3_CalP1_SP0_GP9_17_Xo2(M3_CalP1_SP0_GP9_17_NotA, vdd, M3_CalP1_SP0_GP9_17_line2);
nand2 M3_CalP1_SP0_GP9_17_Xo3(M3_CalP1_SP0_GP9_17_NotB, Xbus_8, M3_CalP1_SP0_GP9_17_line3);
nand2 M3_CalP1_SP0_GP9_17_Xo4(M3_CalP1_SP0_GP9_17_line2, M3_CalP1_SP0_GP9_17_line3, M3_CalP1_Propbus_8);
or2 M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_0(M3_CalP1_Genbus_0, M3_CalP1_Propbus_0, M3_CalP1_LocalC1_0);
and2 M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_1_Ao2_0(M3_CalP1_Propbus_1, M3_CalP1_Genbus_0, M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_1_line0);
or2 M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_1_Ao2_1(M3_CalP1_Genbus_1, M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_1_line0, M3_CalP1_LocalC0_1);
and2 M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_2_Ao3a_0(M3_CalP1_Propbus_1, M3_CalP1_Genbus_0, M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_2_line0);
and2 M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_2_Ao3a_1(M3_CalP1_Propbus_1, M3_CalP1_Propbus_0, M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_2_line1);
or3 M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_2_Ao3a_2(M3_CalP1_Genbus_1, M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_2_line0, M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_2_line1, M3_CalP1_LocalC1_1);
and2 M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_3_Ao3a_0(M3_CalP1_Propbus_2, M3_CalP1_Genbus_1, M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_3_line0);
and3 M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_3_Ao3a_1(M3_CalP1_Propbus_2, M3_CalP1_Propbus_1, M3_CalP1_Genbus_0, M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_3_line1);
or3 M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_3_Ao3a_2(M3_CalP1_Genbus_2, M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_3_line0, M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_3_line1, M3_CalP1_LocalC0_2);
and2 M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_4_Ao4a_0(M3_CalP1_Propbus_2, M3_CalP1_Genbus_1, M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_4_line0);
and3 M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_4_Ao4a_1(M3_CalP1_Propbus_2, M3_CalP1_Propbus_1, M3_CalP1_Genbus_0, M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_4_line1);
and3 M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_4_Ao4a_2(M3_CalP1_Propbus_2, M3_CalP1_Propbus_1, M3_CalP1_Propbus_0, M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_4_line2);
or4 M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_4_Ao4a_3(M3_CalP1_Genbus_2, M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_4_line0, M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_4_line1, M3_CalP1_SP1_GLC5_0_GLC4_0_GLC4_4_line2, M3_CalP1_LocalC1_2);
and2 M3_CalP1_SP1_GLC5_0_GLC4_1_Ao4a_0(M3_CalP1_Propbus_3, M3_CalP1_Genbus_2, M3_CalP1_SP1_GLC5_0_GLC4_1_line0);
and3 M3_CalP1_SP1_GLC5_0_GLC4_1_Ao4a_1(M3_CalP1_Propbus_3, M3_CalP1_Propbus_2, M3_CalP1_Genbus_1, M3_CalP1_SP1_GLC5_0_GLC4_1_line1);
and4 M3_CalP1_SP1_GLC5_0_GLC4_1_Ao4a_2(M3_CalP1_Propbus_3, M3_CalP1_Propbus_2, M3_CalP1_Propbus_1, M3_CalP1_Genbus_0, M3_CalP1_SP1_GLC5_0_GLC4_1_line2);
or4 M3_CalP1_SP1_GLC5_0_GLC4_1_Ao4a_3(M3_CalP1_Genbus_3, M3_CalP1_SP1_GLC5_0_GLC4_1_line0, M3_CalP1_SP1_GLC5_0_GLC4_1_line1, M3_CalP1_SP1_GLC5_0_GLC4_1_line2, M3_CalP1_LocalC0_3);
and2 M3_CalP1_SP1_GLC5_0_GLC4_2_Ao5a_0(M3_CalP1_Propbus_3, M3_CalP1_Genbus_2, M3_CalP1_SP1_GLC5_0_GLC4_2_line0);
and3 M3_CalP1_SP1_GLC5_0_GLC4_2_Ao5a_1(M3_CalP1_Propbus_3, M3_CalP1_Propbus_2, M3_CalP1_Genbus_1, M3_CalP1_SP1_GLC5_0_GLC4_2_line1);
and4 M3_CalP1_SP1_GLC5_0_GLC4_2_Ao5a_2(M3_CalP1_Propbus_3, M3_CalP1_Propbus_2, M3_CalP1_Propbus_1, M3_CalP1_Genbus_0, M3_CalP1_SP1_GLC5_0_GLC4_2_line2);
and4 M3_CalP1_SP1_GLC5_0_GLC4_2_Ao5a_3(M3_CalP1_Propbus_3, M3_CalP1_Propbus_2, M3_CalP1_Propbus_1, M3_CalP1_Propbus_0, M3_CalP1_SP1_GLC5_0_GLC4_2_line3);
or5 M3_CalP1_SP1_GLC5_0_GLC4_2_Ao5a_4(M3_CalP1_Genbus_3, M3_CalP1_SP1_GLC5_0_GLC4_2_line0, M3_CalP1_SP1_GLC5_0_GLC4_2_line1, M3_CalP1_SP1_GLC5_0_GLC4_2_line2, M3_CalP1_SP1_GLC5_0_GLC4_2_line3, M3_CalP1_LocalC1_3);
and2 M3_CalP1_SP1_GLC5_1_Ao5a_0(M3_CalP1_Propbus_4, M3_CalP1_Genbus_3, M3_CalP1_SP1_GLC5_1_line0);
and3 M3_CalP1_SP1_GLC5_1_Ao5a_1(M3_CalP1_Propbus_4, M3_CalP1_Propbus_3, M3_CalP1_Genbus_2, M3_CalP1_SP1_GLC5_1_line1);
and4 M3_CalP1_SP1_GLC5_1_Ao5a_2(M3_CalP1_Propbus_4, M3_CalP1_Propbus_3, M3_CalP1_Propbus_2, M3_CalP1_Genbus_1, M3_CalP1_SP1_GLC5_1_line2);
and5 M3_CalP1_SP1_GLC5_1_Ao5a_3(M3_CalP1_Propbus_4, M3_CalP1_Propbus_3, M3_CalP1_Propbus_2, M3_CalP1_Propbus_1, M3_CalP1_Genbus_0, M3_CalP1_SP1_GLC5_1_line3);
or5 M3_CalP1_SP1_GLC5_1_Ao5a_4(M3_CalP1_Genbus_4, M3_CalP1_SP1_GLC5_1_line0, M3_CalP1_SP1_GLC5_1_line1, M3_CalP1_SP1_GLC5_1_line2, M3_CalP1_SP1_GLC5_1_line3, M3_CalP1_LocalC0_4);
and2 M3_CalP1_SP1_GLC5_2_Ao6a_0(M3_CalP1_Propbus_4, M3_CalP1_Genbus_3, M3_CalP1_SP1_GLC5_2_line0);
and3 M3_CalP1_SP1_GLC5_2_Ao6a_1(M3_CalP1_Propbus_4, M3_CalP1_Propbus_3, M3_CalP1_Genbus_2, M3_CalP1_SP1_GLC5_2_line1);
and4 M3_CalP1_SP1_GLC5_2_Ao6a_2(M3_CalP1_Propbus_4, M3_CalP1_Propbus_3, M3_CalP1_Propbus_2, M3_CalP1_Genbus_1, M3_CalP1_SP1_GLC5_2_line2);
and5 M3_CalP1_SP1_GLC5_2_Ao6a_3(M3_CalP1_Propbus_4, M3_CalP1_Propbus_3, M3_CalP1_Propbus_2, M3_CalP1_Propbus_1, M3_CalP1_Genbus_0, M3_CalP1_SP1_GLC5_2_line3);
and5 M3_CalP1_SP1_GLC5_2_Ao6a_4(M3_CalP1_Propbus_4, M3_CalP1_Propbus_3, M3_CalP1_Propbus_2, M3_CalP1_Propbus_1, M3_CalP1_Propbus_0, M3_CalP1_SP1_GLC5_2_line4);
or6 M3_CalP1_SP1_GLC5_2_Ao6a_5(M3_CalP1_Genbus_4, M3_CalP1_SP1_GLC5_2_line0, M3_CalP1_SP1_GLC5_2_line1, M3_CalP1_SP1_GLC5_2_line2, M3_CalP1_SP1_GLC5_2_line3, M3_CalP1_SP1_GLC5_2_line4, M3_CalP1_LocalC1_4);
or2 M3_CalP1_SP2_GLC4_0(M3_CalP1_Genbus_5, M3_CalP1_Propbus_5, M3_CalP1_LocalC1_5);
and2 M3_CalP1_SP2_GLC4_1_Ao2_0(M3_CalP1_Propbus_6, M3_CalP1_Genbus_5, M3_CalP1_SP2_GLC4_1_line0);
or2 M3_CalP1_SP2_GLC4_1_Ao2_1(M3_CalP1_Genbus_6, M3_CalP1_SP2_GLC4_1_line0, M3_CalP1_LocalC0_6);
and2 M3_CalP1_SP2_GLC4_2_Ao3a_0(M3_CalP1_Propbus_6, M3_CalP1_Genbus_5, M3_CalP1_SP2_GLC4_2_line0);
and2 M3_CalP1_SP2_GLC4_2_Ao3a_1(M3_CalP1_Propbus_6, M3_CalP1_Propbus_5, M3_CalP1_SP2_GLC4_2_line1);
or3 M3_CalP1_SP2_GLC4_2_Ao3a_2(M3_CalP1_Genbus_6, M3_CalP1_SP2_GLC4_2_line0, M3_CalP1_SP2_GLC4_2_line1, M3_CalP1_LocalC1_6);
and2 M3_CalP1_SP2_GLC4_3_Ao3a_0(M3_CalP1_Propbus_7, M3_CalP1_Genbus_6, M3_CalP1_SP2_GLC4_3_line0);
and3 M3_CalP1_SP2_GLC4_3_Ao3a_1(M3_CalP1_Propbus_7, M3_CalP1_Propbus_6, M3_CalP1_Genbus_5, M3_CalP1_SP2_GLC4_3_line1);
or3 M3_CalP1_SP2_GLC4_3_Ao3a_2(M3_CalP1_Genbus_7, M3_CalP1_SP2_GLC4_3_line0, M3_CalP1_SP2_GLC4_3_line1, M3_CalP1_LocalC0_7);
and2 M3_CalP1_SP2_GLC4_4_Ao4a_0(M3_CalP1_Propbus_7, M3_CalP1_Genbus_6, M3_CalP1_SP2_GLC4_4_line0);
and3 M3_CalP1_SP2_GLC4_4_Ao4a_1(M3_CalP1_Propbus_7, M3_CalP1_Propbus_6, M3_CalP1_Genbus_5, M3_CalP1_SP2_GLC4_4_line1);
and3 M3_CalP1_SP2_GLC4_4_Ao4a_2(M3_CalP1_Propbus_7, M3_CalP1_Propbus_6, M3_CalP1_Propbus_5, M3_CalP1_SP2_GLC4_4_line2);
or4 M3_CalP1_SP2_GLC4_4_Ao4a_3(M3_CalP1_Genbus_7, M3_CalP1_SP2_GLC4_4_line0, M3_CalP1_SP2_GLC4_4_line1, M3_CalP1_SP2_GLC4_4_line2, M3_CalP1_LocalC1_7);
inv M3_CalP1_SP3_SP9nc0_SP7nc0_Xo0(M3_CalP1_Genbus_0, M3_CalP1_SP3_SP9nc0_SP7nc0_NotA);
inv M3_CalP1_SP3_SP9nc0_SP7nc0_Xo1(M3_CalP1_LocalC0_1, M3_CalP1_SP3_SP9nc0_SP7nc0_NotB);
nand2 M3_CalP1_SP3_SP9nc0_SP7nc0_Xo2(M3_CalP1_SP3_SP9nc0_SP7nc0_NotA, M3_CalP1_LocalC0_1, M3_CalP1_SP3_SP9nc0_SP7nc0_line2);
nand2 M3_CalP1_SP3_SP9nc0_SP7nc0_Xo3(M3_CalP1_SP3_SP9nc0_SP7nc0_NotB, M3_CalP1_Genbus_0, M3_CalP1_SP3_SP9nc0_SP7nc0_line3);
nand2 M3_CalP1_SP3_SP9nc0_SP7nc0_Xo4(M3_CalP1_SP3_SP9nc0_SP7nc0_line2, M3_CalP1_SP3_SP9nc0_SP7nc0_line3, M3_CalP1_SP3_SP9nc0_line0);
inv M3_CalP1_SP3_SP9nc0_SP7nc1_Xo0(M3_CalP1_LocalC0_2, M3_CalP1_SP3_SP9nc0_SP7nc1_NotA);
inv M3_CalP1_SP3_SP9nc0_SP7nc1_Xo1(M3_CalP1_SP3_SP9nc0_line0, M3_CalP1_SP3_SP9nc0_SP7nc1_NotB);
nand2 M3_CalP1_SP3_SP9nc0_SP7nc1_Xo2(M3_CalP1_SP3_SP9nc0_SP7nc1_NotA, M3_CalP1_SP3_SP9nc0_line0, M3_CalP1_SP3_SP9nc0_SP7nc1_line2);
nand2 M3_CalP1_SP3_SP9nc0_SP7nc1_Xo3(M3_CalP1_SP3_SP9nc0_SP7nc1_NotB, M3_CalP1_LocalC0_2, M3_CalP1_SP3_SP9nc0_SP7nc1_line3);
nand2 M3_CalP1_SP3_SP9nc0_SP7nc1_Xo4(M3_CalP1_SP3_SP9nc0_SP7nc1_line2, M3_CalP1_SP3_SP9nc0_SP7nc1_line3, M3_CalP1_SP3_SP9nc0_line1);
inv M3_CalP1_SP3_SP9nc0_SP7nc2_Xo0(M3_CalP1_LocalC0_3, M3_CalP1_SP3_SP9nc0_SP7nc2_NotA);
inv M3_CalP1_SP3_SP9nc0_SP7nc2_Xo1(M3_CalP1_SP3_SP9nc0_line1, M3_CalP1_SP3_SP9nc0_SP7nc2_NotB);
nand2 M3_CalP1_SP3_SP9nc0_SP7nc2_Xo2(M3_CalP1_SP3_SP9nc0_SP7nc2_NotA, M3_CalP1_SP3_SP9nc0_line1, M3_CalP1_SP3_SP9nc0_SP7nc2_line2);
nand2 M3_CalP1_SP3_SP9nc0_SP7nc2_Xo3(M3_CalP1_SP3_SP9nc0_SP7nc2_NotB, M3_CalP1_LocalC0_3, M3_CalP1_SP3_SP9nc0_SP7nc2_line3);
nand2 M3_CalP1_SP3_SP9nc0_SP7nc2_Xo4(M3_CalP1_SP3_SP9nc0_SP7nc2_line2, M3_CalP1_SP3_SP9nc0_SP7nc2_line3, M3_CalP1_SP3_SP9nc0_line2);
inv M3_CalP1_SP3_SP9nc0_SP7nc3_Xo0(M3_CalP1_Propbus_0, M3_CalP1_SP3_SP9nc0_SP7nc3_NotA);
inv M3_CalP1_SP3_SP9nc0_SP7nc3_Xo1(M3_CalP1_SP3_SP9nc0_line2, M3_CalP1_SP3_SP9nc0_SP7nc3_NotB);
nand2 M3_CalP1_SP3_SP9nc0_SP7nc3_Xo2(M3_CalP1_SP3_SP9nc0_SP7nc3_NotA, M3_CalP1_SP3_SP9nc0_line2, M3_CalP1_SP3_SP9nc0_SP7nc3_line2);
nand2 M3_CalP1_SP3_SP9nc0_SP7nc3_Xo3(M3_CalP1_SP3_SP9nc0_SP7nc3_NotB, M3_CalP1_Propbus_0, M3_CalP1_SP3_SP9nc0_SP7nc3_line3);
nand2 M3_CalP1_SP3_SP9nc0_SP7nc3_Xo4(M3_CalP1_SP3_SP9nc0_SP7nc3_line2, M3_CalP1_SP3_SP9nc0_SP7nc3_line3, M3_CalP1_SP3_SP9nc0_line3);
inv M3_CalP1_SP3_SP9nc0_SP7nc4_Xo0(M3_CalP1_Propbus_1, M3_CalP1_SP3_SP9nc0_SP7nc4_NotA);
inv M3_CalP1_SP3_SP9nc0_SP7nc4_Xo1(M3_CalP1_SP3_SP9nc0_line3, M3_CalP1_SP3_SP9nc0_SP7nc4_NotB);
nand2 M3_CalP1_SP3_SP9nc0_SP7nc4_Xo2(M3_CalP1_SP3_SP9nc0_SP7nc4_NotA, M3_CalP1_SP3_SP9nc0_line3, M3_CalP1_SP3_SP9nc0_SP7nc4_line2);
nand2 M3_CalP1_SP3_SP9nc0_SP7nc4_Xo3(M3_CalP1_SP3_SP9nc0_SP7nc4_NotB, M3_CalP1_Propbus_1, M3_CalP1_SP3_SP9nc0_SP7nc4_line3);
nand2 M3_CalP1_SP3_SP9nc0_SP7nc4_Xo4(M3_CalP1_SP3_SP9nc0_SP7nc4_line2, M3_CalP1_SP3_SP9nc0_SP7nc4_line3, M3_CalP1_SP3_SP9nc0_line4);
inv M3_CalP1_SP3_SP9nc0_SP7nc5_Xo0(M3_CalP1_Propbus_2, M3_CalP1_SP3_SP9nc0_SP7nc5_NotA);
inv M3_CalP1_SP3_SP9nc0_SP7nc5_Xo1(M3_CalP1_SP3_SP9nc0_line4, M3_CalP1_SP3_SP9nc0_SP7nc5_NotB);
nand2 M3_CalP1_SP3_SP9nc0_SP7nc5_Xo2(M3_CalP1_SP3_SP9nc0_SP7nc5_NotA, M3_CalP1_SP3_SP9nc0_line4, M3_CalP1_SP3_SP9nc0_SP7nc5_line2);
nand2 M3_CalP1_SP3_SP9nc0_SP7nc5_Xo3(M3_CalP1_SP3_SP9nc0_SP7nc5_NotB, M3_CalP1_Propbus_2, M3_CalP1_SP3_SP9nc0_SP7nc5_line3);
nand2 M3_CalP1_SP3_SP9nc0_SP7nc5_Xo4(M3_CalP1_SP3_SP9nc0_SP7nc5_line2, M3_CalP1_SP3_SP9nc0_SP7nc5_line3, M3_CalP1_SP3_line0);
inv M3_CalP1_SP3_SP9nc1_Xo0(M3_CalP1_Propbus_3, M3_CalP1_SP3_SP9nc1_NotA);
inv M3_CalP1_SP3_SP9nc1_Xo1(M3_CalP1_SP3_line0, M3_CalP1_SP3_SP9nc1_NotB);
nand2 M3_CalP1_SP3_SP9nc1_Xo2(M3_CalP1_SP3_SP9nc1_NotA, M3_CalP1_SP3_line0, M3_CalP1_SP3_SP9nc1_line2);
nand2 M3_CalP1_SP3_SP9nc1_Xo3(M3_CalP1_SP3_SP9nc1_NotB, M3_CalP1_Propbus_3, M3_CalP1_SP3_SP9nc1_line3);
nand2 M3_CalP1_SP3_SP9nc1_Xo4(M3_CalP1_SP3_SP9nc1_line2, M3_CalP1_SP3_SP9nc1_line3, M3_CalP1_SP3_line1);
inv M3_CalP1_SP3_SP9nc2_Xo0(M3_CalP1_Propbus_4, M3_CalP1_SP3_SP9nc2_NotA);
inv M3_CalP1_SP3_SP9nc2_Xo1(M3_CalP1_SP3_line1, M3_CalP1_SP3_SP9nc2_NotB);
nand2 M3_CalP1_SP3_SP9nc2_Xo2(M3_CalP1_SP3_SP9nc2_NotA, M3_CalP1_SP3_line1, M3_CalP1_SP3_SP9nc2_line2);
nand2 M3_CalP1_SP3_SP9nc2_Xo3(M3_CalP1_SP3_SP9nc2_NotB, M3_CalP1_Propbus_4, M3_CalP1_SP3_SP9nc2_line3);
nand2 M3_CalP1_SP3_SP9nc2_Xo4(M3_CalP1_SP3_SP9nc2_line2, M3_CalP1_SP3_SP9nc2_line3, M3_CalP1_ParLo0);
inv M3_CalP1_SP4_SP9nc0_SP7c0(M3_CalP1_Propbus_2, M3_CalP1_SP4_SP9nc0_NewInbus_6);
inv M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_Xo0(M3_CalP1_LocalC1_0, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_NotA);
inv M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_Xo1(M3_CalP1_LocalC1_1, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_NotB);
nand2 M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_Xo2(M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_NotA, M3_CalP1_LocalC1_1, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_line2);
nand2 M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_Xo3(M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_NotB, M3_CalP1_LocalC1_0, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_line3);
nand2 M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_Xo4(M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_line2, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_line3, M3_CalP1_SP4_SP9nc0_SP7c2_line0);
inv M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_Xo0(M3_CalP1_LocalC1_2, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_NotA);
inv M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_Xo1(M3_CalP1_SP4_SP9nc0_SP7c2_line0, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_NotB);
nand2 M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_Xo2(M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_NotA, M3_CalP1_SP4_SP9nc0_SP7c2_line0, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_line2);
nand2 M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_Xo3(M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_NotB, M3_CalP1_LocalC1_2, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_line3);
nand2 M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_Xo4(M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_line2, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_line3, M3_CalP1_SP4_SP9nc0_SP7c2_line1);
inv M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_Xo0(M3_CalP1_LocalC1_3, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_NotA);
inv M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_Xo1(M3_CalP1_SP4_SP9nc0_SP7c2_line1, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_NotB);
nand2 M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_Xo2(M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_NotA, M3_CalP1_SP4_SP9nc0_SP7c2_line1, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_line2);
nand2 M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_Xo3(M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_NotB, M3_CalP1_LocalC1_3, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_line3);
nand2 M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_Xo4(M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_line2, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_line3, M3_CalP1_SP4_SP9nc0_SP7c2_line2);
inv M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_Xo0(M3_CalP1_Propbus_0, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_NotA);
inv M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_Xo1(M3_CalP1_SP4_SP9nc0_SP7c2_line2, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_NotB);
nand2 M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_Xo2(M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_NotA, M3_CalP1_SP4_SP9nc0_SP7c2_line2, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_line2);
nand2 M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_Xo3(M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_NotB, M3_CalP1_Propbus_0, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_line3);
nand2 M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_Xo4(M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_line2, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_line3, M3_CalP1_SP4_SP9nc0_SP7c2_line3);
inv M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_Xo0(M3_CalP1_Propbus_1, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_NotA);
inv M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_Xo1(M3_CalP1_SP4_SP9nc0_SP7c2_line3, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_NotB);
nand2 M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_Xo2(M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_NotA, M3_CalP1_SP4_SP9nc0_SP7c2_line3, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_line2);
nand2 M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_Xo3(M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_NotB, M3_CalP1_Propbus_1, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_line3);
nand2 M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_Xo4(M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_line2, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_line3, M3_CalP1_SP4_SP9nc0_SP7c2_line4);
inv M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_Xo0(M3_CalP1_SP4_SP9nc0_NewInbus_6, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_NotA);
inv M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_Xo1(M3_CalP1_SP4_SP9nc0_SP7c2_line4, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_NotB);
nand2 M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_Xo2(M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_NotA, M3_CalP1_SP4_SP9nc0_SP7c2_line4, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_line2);
nand2 M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_Xo3(M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_NotB, M3_CalP1_SP4_SP9nc0_NewInbus_6, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_line3);
nand2 M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_Xo4(M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_line2, M3_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_line3, M3_CalP1_SP4_line0);
inv M3_CalP1_SP4_SP9nc1_Xo0(M3_CalP1_Propbus_3, M3_CalP1_SP4_SP9nc1_NotA);
inv M3_CalP1_SP4_SP9nc1_Xo1(M3_CalP1_SP4_line0, M3_CalP1_SP4_SP9nc1_NotB);
nand2 M3_CalP1_SP4_SP9nc1_Xo2(M3_CalP1_SP4_SP9nc1_NotA, M3_CalP1_SP4_line0, M3_CalP1_SP4_SP9nc1_line2);
nand2 M3_CalP1_SP4_SP9nc1_Xo3(M3_CalP1_SP4_SP9nc1_NotB, M3_CalP1_Propbus_3, M3_CalP1_SP4_SP9nc1_line3);
nand2 M3_CalP1_SP4_SP9nc1_Xo4(M3_CalP1_SP4_SP9nc1_line2, M3_CalP1_SP4_SP9nc1_line3, M3_CalP1_SP4_line1);
inv M3_CalP1_SP4_SP9nc2_Xo0(M3_CalP1_Propbus_4, M3_CalP1_SP4_SP9nc2_NotA);
inv M3_CalP1_SP4_SP9nc2_Xo1(M3_CalP1_SP4_line1, M3_CalP1_SP4_SP9nc2_NotB);
nand2 M3_CalP1_SP4_SP9nc2_Xo2(M3_CalP1_SP4_SP9nc2_NotA, M3_CalP1_SP4_line1, M3_CalP1_SP4_SP9nc2_line2);
nand2 M3_CalP1_SP4_SP9nc2_Xo3(M3_CalP1_SP4_SP9nc2_NotB, M3_CalP1_Propbus_4, M3_CalP1_SP4_SP9nc2_line3);
nand2 M3_CalP1_SP4_SP9nc2_Xo4(M3_CalP1_SP4_SP9nc2_line2, M3_CalP1_SP4_SP9nc2_line3, M3_CalP1_ParLo1);
inv M3_CalP1_SP5_SP7nc0_Xo0(M3_CalP1_Genbus_5, M3_CalP1_SP5_SP7nc0_NotA);
inv M3_CalP1_SP5_SP7nc0_Xo1(M3_CalP1_LocalC0_6, M3_CalP1_SP5_SP7nc0_NotB);
nand2 M3_CalP1_SP5_SP7nc0_Xo2(M3_CalP1_SP5_SP7nc0_NotA, M3_CalP1_LocalC0_6, M3_CalP1_SP5_SP7nc0_line2);
nand2 M3_CalP1_SP5_SP7nc0_Xo3(M3_CalP1_SP5_SP7nc0_NotB, M3_CalP1_Genbus_5, M3_CalP1_SP5_SP7nc0_line3);
nand2 M3_CalP1_SP5_SP7nc0_Xo4(M3_CalP1_SP5_SP7nc0_line2, M3_CalP1_SP5_SP7nc0_line3, M3_CalP1_SP5_line0);
inv M3_CalP1_SP5_SP7nc1_Xo0(M3_CalP1_LocalC0_7, M3_CalP1_SP5_SP7nc1_NotA);
inv M3_CalP1_SP5_SP7nc1_Xo1(M3_CalP1_SP5_line0, M3_CalP1_SP5_SP7nc1_NotB);
nand2 M3_CalP1_SP5_SP7nc1_Xo2(M3_CalP1_SP5_SP7nc1_NotA, M3_CalP1_SP5_line0, M3_CalP1_SP5_SP7nc1_line2);
nand2 M3_CalP1_SP5_SP7nc1_Xo3(M3_CalP1_SP5_SP7nc1_NotB, M3_CalP1_LocalC0_7, M3_CalP1_SP5_SP7nc1_line3);
nand2 M3_CalP1_SP5_SP7nc1_Xo4(M3_CalP1_SP5_SP7nc1_line2, M3_CalP1_SP5_SP7nc1_line3, M3_CalP1_SP5_line1);
inv M3_CalP1_SP5_SP7nc2_Xo0(M3_CalP1_Propbus_5, M3_CalP1_SP5_SP7nc2_NotA);
inv M3_CalP1_SP5_SP7nc2_Xo1(M3_CalP1_SP5_line1, M3_CalP1_SP5_SP7nc2_NotB);
nand2 M3_CalP1_SP5_SP7nc2_Xo2(M3_CalP1_SP5_SP7nc2_NotA, M3_CalP1_SP5_line1, M3_CalP1_SP5_SP7nc2_line2);
nand2 M3_CalP1_SP5_SP7nc2_Xo3(M3_CalP1_SP5_SP7nc2_NotB, M3_CalP1_Propbus_5, M3_CalP1_SP5_SP7nc2_line3);
nand2 M3_CalP1_SP5_SP7nc2_Xo4(M3_CalP1_SP5_SP7nc2_line2, M3_CalP1_SP5_SP7nc2_line3, M3_CalP1_SP5_line2);
inv M3_CalP1_SP5_SP7nc3_Xo0(M3_CalP1_Propbus_6, M3_CalP1_SP5_SP7nc3_NotA);
inv M3_CalP1_SP5_SP7nc3_Xo1(M3_CalP1_SP5_line2, M3_CalP1_SP5_SP7nc3_NotB);
nand2 M3_CalP1_SP5_SP7nc3_Xo2(M3_CalP1_SP5_SP7nc3_NotA, M3_CalP1_SP5_line2, M3_CalP1_SP5_SP7nc3_line2);
nand2 M3_CalP1_SP5_SP7nc3_Xo3(M3_CalP1_SP5_SP7nc3_NotB, M3_CalP1_Propbus_6, M3_CalP1_SP5_SP7nc3_line3);
nand2 M3_CalP1_SP5_SP7nc3_Xo4(M3_CalP1_SP5_SP7nc3_line2, M3_CalP1_SP5_SP7nc3_line3, M3_CalP1_SP5_line3);
inv M3_CalP1_SP5_SP7nc4_Xo0(M3_CalP1_Propbus_7, M3_CalP1_SP5_SP7nc4_NotA);
inv M3_CalP1_SP5_SP7nc4_Xo1(M3_CalP1_SP5_line3, M3_CalP1_SP5_SP7nc4_NotB);
nand2 M3_CalP1_SP5_SP7nc4_Xo2(M3_CalP1_SP5_SP7nc4_NotA, M3_CalP1_SP5_line3, M3_CalP1_SP5_SP7nc4_line2);
nand2 M3_CalP1_SP5_SP7nc4_Xo3(M3_CalP1_SP5_SP7nc4_NotB, M3_CalP1_Propbus_7, M3_CalP1_SP5_SP7nc4_line3);
nand2 M3_CalP1_SP5_SP7nc4_Xo4(M3_CalP1_SP5_SP7nc4_line2, M3_CalP1_SP5_SP7nc4_line3, M3_CalP1_SP5_line4);
inv M3_CalP1_SP5_SP7nc5_Xo0(M3_CalP1_Propbus_8, M3_CalP1_SP5_SP7nc5_NotA);
inv M3_CalP1_SP5_SP7nc5_Xo1(M3_CalP1_SP5_line4, M3_CalP1_SP5_SP7nc5_NotB);
nand2 M3_CalP1_SP5_SP7nc5_Xo2(M3_CalP1_SP5_SP7nc5_NotA, M3_CalP1_SP5_line4, M3_CalP1_SP5_SP7nc5_line2);
nand2 M3_CalP1_SP5_SP7nc5_Xo3(M3_CalP1_SP5_SP7nc5_NotB, M3_CalP1_Propbus_8, M3_CalP1_SP5_SP7nc5_line3);
nand2 M3_CalP1_SP5_SP7nc5_Xo4(M3_CalP1_SP5_SP7nc5_line2, M3_CalP1_SP5_SP7nc5_line3, M3_CalP1_ParHi0);
inv M3_CalP1_SP6_SP7c0(M3_CalP1_Propbus_8, M3_CalP1_SP6_NewInbus_6);
inv M3_CalP1_SP6_SP7c2_SP7nc0_Xo0(M3_CalP1_LocalC1_5, M3_CalP1_SP6_SP7c2_SP7nc0_NotA);
inv M3_CalP1_SP6_SP7c2_SP7nc0_Xo1(M3_CalP1_LocalC1_6, M3_CalP1_SP6_SP7c2_SP7nc0_NotB);
nand2 M3_CalP1_SP6_SP7c2_SP7nc0_Xo2(M3_CalP1_SP6_SP7c2_SP7nc0_NotA, M3_CalP1_LocalC1_6, M3_CalP1_SP6_SP7c2_SP7nc0_line2);
nand2 M3_CalP1_SP6_SP7c2_SP7nc0_Xo3(M3_CalP1_SP6_SP7c2_SP7nc0_NotB, M3_CalP1_LocalC1_5, M3_CalP1_SP6_SP7c2_SP7nc0_line3);
nand2 M3_CalP1_SP6_SP7c2_SP7nc0_Xo4(M3_CalP1_SP6_SP7c2_SP7nc0_line2, M3_CalP1_SP6_SP7c2_SP7nc0_line3, M3_CalP1_SP6_SP7c2_line0);
inv M3_CalP1_SP6_SP7c2_SP7nc1_Xo0(M3_CalP1_LocalC1_7, M3_CalP1_SP6_SP7c2_SP7nc1_NotA);
inv M3_CalP1_SP6_SP7c2_SP7nc1_Xo1(M3_CalP1_SP6_SP7c2_line0, M3_CalP1_SP6_SP7c2_SP7nc1_NotB);
nand2 M3_CalP1_SP6_SP7c2_SP7nc1_Xo2(M3_CalP1_SP6_SP7c2_SP7nc1_NotA, M3_CalP1_SP6_SP7c2_line0, M3_CalP1_SP6_SP7c2_SP7nc1_line2);
nand2 M3_CalP1_SP6_SP7c2_SP7nc1_Xo3(M3_CalP1_SP6_SP7c2_SP7nc1_NotB, M3_CalP1_LocalC1_7, M3_CalP1_SP6_SP7c2_SP7nc1_line3);
nand2 M3_CalP1_SP6_SP7c2_SP7nc1_Xo4(M3_CalP1_SP6_SP7c2_SP7nc1_line2, M3_CalP1_SP6_SP7c2_SP7nc1_line3, M3_CalP1_SP6_SP7c2_line1);
inv M3_CalP1_SP6_SP7c2_SP7nc2_Xo0(M3_CalP1_Propbus_5, M3_CalP1_SP6_SP7c2_SP7nc2_NotA);
inv M3_CalP1_SP6_SP7c2_SP7nc2_Xo1(M3_CalP1_SP6_SP7c2_line1, M3_CalP1_SP6_SP7c2_SP7nc2_NotB);
nand2 M3_CalP1_SP6_SP7c2_SP7nc2_Xo2(M3_CalP1_SP6_SP7c2_SP7nc2_NotA, M3_CalP1_SP6_SP7c2_line1, M3_CalP1_SP6_SP7c2_SP7nc2_line2);
nand2 M3_CalP1_SP6_SP7c2_SP7nc2_Xo3(M3_CalP1_SP6_SP7c2_SP7nc2_NotB, M3_CalP1_Propbus_5, M3_CalP1_SP6_SP7c2_SP7nc2_line3);
nand2 M3_CalP1_SP6_SP7c2_SP7nc2_Xo4(M3_CalP1_SP6_SP7c2_SP7nc2_line2, M3_CalP1_SP6_SP7c2_SP7nc2_line3, M3_CalP1_SP6_SP7c2_line2);
inv M3_CalP1_SP6_SP7c2_SP7nc3_Xo0(M3_CalP1_Propbus_6, M3_CalP1_SP6_SP7c2_SP7nc3_NotA);
inv M3_CalP1_SP6_SP7c2_SP7nc3_Xo1(M3_CalP1_SP6_SP7c2_line2, M3_CalP1_SP6_SP7c2_SP7nc3_NotB);
nand2 M3_CalP1_SP6_SP7c2_SP7nc3_Xo2(M3_CalP1_SP6_SP7c2_SP7nc3_NotA, M3_CalP1_SP6_SP7c2_line2, M3_CalP1_SP6_SP7c2_SP7nc3_line2);
nand2 M3_CalP1_SP6_SP7c2_SP7nc3_Xo3(M3_CalP1_SP6_SP7c2_SP7nc3_NotB, M3_CalP1_Propbus_6, M3_CalP1_SP6_SP7c2_SP7nc3_line3);
nand2 M3_CalP1_SP6_SP7c2_SP7nc3_Xo4(M3_CalP1_SP6_SP7c2_SP7nc3_line2, M3_CalP1_SP6_SP7c2_SP7nc3_line3, M3_CalP1_SP6_SP7c2_line3);
inv M3_CalP1_SP6_SP7c2_SP7nc4_Xo0(M3_CalP1_Propbus_7, M3_CalP1_SP6_SP7c2_SP7nc4_NotA);
inv M3_CalP1_SP6_SP7c2_SP7nc4_Xo1(M3_CalP1_SP6_SP7c2_line3, M3_CalP1_SP6_SP7c2_SP7nc4_NotB);
nand2 M3_CalP1_SP6_SP7c2_SP7nc4_Xo2(M3_CalP1_SP6_SP7c2_SP7nc4_NotA, M3_CalP1_SP6_SP7c2_line3, M3_CalP1_SP6_SP7c2_SP7nc4_line2);
nand2 M3_CalP1_SP6_SP7c2_SP7nc4_Xo3(M3_CalP1_SP6_SP7c2_SP7nc4_NotB, M3_CalP1_Propbus_7, M3_CalP1_SP6_SP7c2_SP7nc4_line3);
nand2 M3_CalP1_SP6_SP7c2_SP7nc4_Xo4(M3_CalP1_SP6_SP7c2_SP7nc4_line2, M3_CalP1_SP6_SP7c2_SP7nc4_line3, M3_CalP1_SP6_SP7c2_line4);
inv M3_CalP1_SP6_SP7c2_SP7nc5_Xo0(M3_CalP1_SP6_NewInbus_6, M3_CalP1_SP6_SP7c2_SP7nc5_NotA);
inv M3_CalP1_SP6_SP7c2_SP7nc5_Xo1(M3_CalP1_SP6_SP7c2_line4, M3_CalP1_SP6_SP7c2_SP7nc5_NotB);
nand2 M3_CalP1_SP6_SP7c2_SP7nc5_Xo2(M3_CalP1_SP6_SP7c2_SP7nc5_NotA, M3_CalP1_SP6_SP7c2_line4, M3_CalP1_SP6_SP7c2_SP7nc5_line2);
nand2 M3_CalP1_SP6_SP7c2_SP7nc5_Xo3(M3_CalP1_SP6_SP7c2_SP7nc5_NotB, M3_CalP1_SP6_NewInbus_6, M3_CalP1_SP6_SP7c2_SP7nc5_line3);
nand2 M3_CalP1_SP6_SP7c2_SP7nc5_Xo4(M3_CalP1_SP6_SP7c2_SP7nc5_line2, M3_CalP1_SP6_SP7c2_SP7nc5_line3, M3_CalP1_ParHi1);
inv M3_CalP1_SP7_Mux2_0(in2174, M3_CalP1_SP7_Not_ContIn);
and2 M3_CalP1_SP7_Mux2_1(M3_CalP1_ParLo0, M3_CalP1_SP7_Not_ContIn, M3_CalP1_SP7_line1);
and2 M3_CalP1_SP7_Mux2_2(M3_CalP1_ParLo1, in2174, M3_CalP1_SP7_line2);
or2 M3_CalP1_SP7_Mux2_3(M3_CalP1_SP7_line1, M3_CalP1_SP7_line2, M3_CalP1_ParLo);
inv M3_CalP1_SP8_Mux2_0(M3_CalP1_LocalC0_4, M3_CalP1_SP8_Not_ContIn);
and2 M3_CalP1_SP8_Mux2_1(M3_CalP1_ParHi0, M3_CalP1_SP8_Not_ContIn, M3_CalP1_SP8_line1);
and2 M3_CalP1_SP8_Mux2_2(M3_CalP1_ParHi1, M3_CalP1_LocalC0_4, M3_CalP1_SP8_line2);
or2 M3_CalP1_SP8_Mux2_3(M3_CalP1_SP8_line1, M3_CalP1_SP8_line2, M3_CalP1_ParHiCin0);
inv M3_CalP1_SP9_Mux2_0(M3_CalP1_LocalC1_4, M3_CalP1_SP9_Not_ContIn);
and2 M3_CalP1_SP9_Mux2_1(M3_CalP1_ParHi0, M3_CalP1_SP9_Not_ContIn, M3_CalP1_SP9_line1);
and2 M3_CalP1_SP9_Mux2_2(M3_CalP1_ParHi1, M3_CalP1_LocalC1_4, M3_CalP1_SP9_line2);
or2 M3_CalP1_SP9_Mux2_3(M3_CalP1_SP9_line1, M3_CalP1_SP9_line2, M3_CalP1_ParHiCin1);
inv M3_CalP1_SP10_Mux2_0(in2174, M3_CalP1_SP10_Not_ContIn);
and2 M3_CalP1_SP10_Mux2_1(M3_CalP1_ParHiCin0, M3_CalP1_SP10_Not_ContIn, M3_CalP1_SP10_line1);
and2 M3_CalP1_SP10_Mux2_2(M3_CalP1_ParHiCin1, in2174, M3_CalP1_SP10_line2);
or2 M3_CalP1_SP10_Mux2_3(M3_CalP1_SP10_line1, M3_CalP1_SP10_line2, M3_CalP1_ParHi);
inv M3_CalP1_SP11_Xo0(M3_CalP1_ParLo, M3_CalP1_SP11_NotA);
inv M3_CalP1_SP11_Xo1(M3_CalP1_ParHi, M3_CalP1_SP11_NotB);
nand2 M3_CalP1_SP11_Xo2(M3_CalP1_SP11_NotA, M3_CalP1_ParHi, M3_CalP1_SP11_line2);
nand2 M3_CalP1_SP11_Xo3(M3_CalP1_SP11_NotB, M3_CalP1_ParLo, M3_CalP1_SP11_line3);
nand2 M3_CalP1_SP11_Xo4(M3_CalP1_SP11_line2, M3_CalP1_SP11_line3, M3_SumPar);
inv M3_CalP2_M2M4_0(M3_LogicPar, M3_CalP2_NotLogicPar);
inv M3_CalP2_M2M4_1(M3_SumPar, M3_CalP2_NotSumPar);
inv M3_CalP2_M2M4_2_Mux2_0(in4091, M3_CalP2_M2M4_2_Not_ContIn);
and2 M3_CalP2_M2M4_2_Mux2_1(M3_CalP2_NotLogicPar, M3_CalP2_M2M4_2_Not_ContIn, M3_CalP2_M2M4_2_line1);
and2 M3_CalP2_M2M4_2_Mux2_2(M3_CalP2_NotSumPar, in4091, M3_CalP2_M2M4_2_line2);
or2 M3_CalP2_M2M4_2_Mux2_3(M3_CalP2_M2M4_2_line1, M3_CalP2_M2M4_2_line2, M3_CalP2_line0);
inv M3_CalP2_M2M4_3_Mux2_0(in4092, M3_CalP2_M2M4_3_Not_ContIn);
and2 M3_CalP2_M2M4_3_Mux2_1(M3_CalP2_line0, M3_CalP2_M2M4_3_Not_ContIn, M3_CalP2_M2M4_3_line1);
and2 M3_CalP2_M2M4_3_Mux2_2(in94, in4092, M3_CalP2_M2M4_3_line2);
or2 M3_CalP2_M2M4_3_Mux2_3(M3_CalP2_M2M4_3_line1, M3_CalP2_M2M4_3_line2, Not_SumLogicParX);
inv M3_CalP2_M2M4_4_Mux4_0(in4092, M3_CalP2_M2M4_4_Not_ContLo);
inv M3_CalP2_M2M4_4_Mux4_1(in4091, M3_CalP2_M2M4_4_Not_ContHi);
and3 M3_CalP2_M2M4_4_Mux4_2(M3_LogicPar, M3_CalP2_M2M4_4_Not_ContHi, M3_CalP2_M2M4_4_Not_ContLo, M3_CalP2_M2M4_4_line2);
and3 M3_CalP2_M2M4_4_Mux4_3(in120, M3_CalP2_M2M4_4_Not_ContHi, in4092, M3_CalP2_M2M4_4_line3);
and3 M3_CalP2_M2M4_4_Mux4_4(M3_SumPar, in4091, M3_CalP2_M2M4_4_Not_ContLo, M3_CalP2_M2M4_4_line4);
and3 M3_CalP2_M2M4_4_Mux4_5(vdd, in4091, in4092, M3_CalP2_M2M4_4_line5);
or4 M3_CalP2_M2M4_4_Mux4_6(M3_CalP2_M2M4_4_line2, M3_CalP2_M2M4_4_line3, M3_CalP2_M2M4_4_line4, M3_CalP2_M2M4_4_line5, out843);
inv M4_CalP0_LP0_CL0_LB0_Mux2_0(in281, M4_CalP0_LP0_CL0_LB0_Not_ContIn);
and2 M4_CalP0_LP0_CL0_LB0_Mux2_1(in254, M4_CalP0_LP0_CL0_LB0_Not_ContIn, M4_CalP0_LP0_CL0_LB0_line1);
and2 M4_CalP0_LP0_CL0_LB0_Mux2_2(in242, in281, M4_CalP0_LP0_CL0_LB0_line2);
or2 M4_CalP0_LP0_CL0_LB0_Mux2_3(M4_CalP0_LP0_CL0_LB0_line1, M4_CalP0_LP0_CL0_LB0_line2, M4_CalP0_LP0_CL0_line0);
inv M4_CalP0_LP0_CL0_LB1_Mux2_0(in281, M4_CalP0_LP0_CL0_LB1_Not_ContIn);
and2 M4_CalP0_LP0_CL0_LB1_Mux2_1(in251, M4_CalP0_LP0_CL0_LB1_Not_ContIn, M4_CalP0_LP0_CL0_LB1_line1);
and2 M4_CalP0_LP0_CL0_LB1_Mux2_2(in248, in281, M4_CalP0_LP0_CL0_LB1_line2);
or2 M4_CalP0_LP0_CL0_LB1_Mux2_3(M4_CalP0_LP0_CL0_LB1_line1, M4_CalP0_LP0_CL0_LB1_line2, M4_CalP0_LP0_CL0_line1);
or2 M4_CalP0_LP0_CL0_LB2(in374, M4_CalP0_LP0_CL0_line0, M4_CalP0_LP0_CL0_line2);
nand2 M4_CalP0_LP0_CL0_LB3(in374, M4_CalP0_LP0_CL0_line1, M4_CalP0_LP0_CL0_line3);
and2 M4_CalP0_LP0_CL0_LB4(M4_CalP0_LP0_CL0_line2, M4_CalP0_LP0_CL0_line3, M4_CalP0_LogicOut_0);
inv M4_CalP0_LP0_CL1_LB0_Mux2_0(in273, M4_CalP0_LP0_CL1_LB0_Not_ContIn);
and2 M4_CalP0_LP0_CL1_LB0_Mux2_1(in254, M4_CalP0_LP0_CL1_LB0_Not_ContIn, M4_CalP0_LP0_CL1_LB0_line1);
and2 M4_CalP0_LP0_CL1_LB0_Mux2_2(in242, in273, M4_CalP0_LP0_CL1_LB0_line2);
or2 M4_CalP0_LP0_CL1_LB0_Mux2_3(M4_CalP0_LP0_CL1_LB0_line1, M4_CalP0_LP0_CL1_LB0_line2, M4_CalP0_LP0_CL1_line0);
inv M4_CalP0_LP0_CL1_LB1_Mux2_0(in273, M4_CalP0_LP0_CL1_LB1_Not_ContIn);
and2 M4_CalP0_LP0_CL1_LB1_Mux2_1(in251, M4_CalP0_LP0_CL1_LB1_Not_ContIn, M4_CalP0_LP0_CL1_LB1_line1);
and2 M4_CalP0_LP0_CL1_LB1_Mux2_2(in248, in273, M4_CalP0_LP0_CL1_LB1_line2);
or2 M4_CalP0_LP0_CL1_LB1_Mux2_3(M4_CalP0_LP0_CL1_LB1_line1, M4_CalP0_LP0_CL1_LB1_line2, M4_CalP0_LP0_CL1_line1);
or2 M4_CalP0_LP0_CL1_LB2(in411, M4_CalP0_LP0_CL1_line0, M4_CalP0_LP0_CL1_line2);
nand2 M4_CalP0_LP0_CL1_LB3(in411, M4_CalP0_LP0_CL1_line1, M4_CalP0_LP0_CL1_line3);
and2 M4_CalP0_LP0_CL1_LB4(M4_CalP0_LP0_CL1_line2, M4_CalP0_LP0_CL1_line3, M4_CalP0_LogicOut_1);
inv M4_CalP0_LP0_CL2_LB0_Mux2_0(in265, M4_CalP0_LP0_CL2_LB0_Not_ContIn);
and2 M4_CalP0_LP0_CL2_LB0_Mux2_1(in254, M4_CalP0_LP0_CL2_LB0_Not_ContIn, M4_CalP0_LP0_CL2_LB0_line1);
and2 M4_CalP0_LP0_CL2_LB0_Mux2_2(in242, in265, M4_CalP0_LP0_CL2_LB0_line2);
or2 M4_CalP0_LP0_CL2_LB0_Mux2_3(M4_CalP0_LP0_CL2_LB0_line1, M4_CalP0_LP0_CL2_LB0_line2, M4_CalP0_LP0_CL2_line0);
inv M4_CalP0_LP0_CL2_LB1_Mux2_0(in265, M4_CalP0_LP0_CL2_LB1_Not_ContIn);
and2 M4_CalP0_LP0_CL2_LB1_Mux2_1(in251, M4_CalP0_LP0_CL2_LB1_Not_ContIn, M4_CalP0_LP0_CL2_LB1_line1);
and2 M4_CalP0_LP0_CL2_LB1_Mux2_2(in248, in265, M4_CalP0_LP0_CL2_LB1_line2);
or2 M4_CalP0_LP0_CL2_LB1_Mux2_3(M4_CalP0_LP0_CL2_LB1_line1, M4_CalP0_LP0_CL2_LB1_line2, M4_CalP0_LP0_CL2_line1);
or2 M4_CalP0_LP0_CL2_LB2(in400, M4_CalP0_LP0_CL2_line0, M4_CalP0_LP0_CL2_line2);
nand2 M4_CalP0_LP0_CL2_LB3(in400, M4_CalP0_LP0_CL2_line1, M4_CalP0_LP0_CL2_line3);
and2 M4_CalP0_LP0_CL2_LB4(M4_CalP0_LP0_CL2_line2, M4_CalP0_LP0_CL2_line3, M4_CalP0_LogicOut_2);
inv M4_CalP0_LP0_CL3_LB0_Mux2_0(in257, M4_CalP0_LP0_CL3_LB0_Not_ContIn);
and2 M4_CalP0_LP0_CL3_LB0_Mux2_1(in254, M4_CalP0_LP0_CL3_LB0_Not_ContIn, M4_CalP0_LP0_CL3_LB0_line1);
and2 M4_CalP0_LP0_CL3_LB0_Mux2_2(in242, in257, M4_CalP0_LP0_CL3_LB0_line2);
or2 M4_CalP0_LP0_CL3_LB0_Mux2_3(M4_CalP0_LP0_CL3_LB0_line1, M4_CalP0_LP0_CL3_LB0_line2, M4_CalP0_LP0_CL3_line0);
inv M4_CalP0_LP0_CL3_LB1_Mux2_0(in257, M4_CalP0_LP0_CL3_LB1_Not_ContIn);
and2 M4_CalP0_LP0_CL3_LB1_Mux2_1(in251, M4_CalP0_LP0_CL3_LB1_Not_ContIn, M4_CalP0_LP0_CL3_LB1_line1);
and2 M4_CalP0_LP0_CL3_LB1_Mux2_2(in248, in257, M4_CalP0_LP0_CL3_LB1_line2);
or2 M4_CalP0_LP0_CL3_LB1_Mux2_3(M4_CalP0_LP0_CL3_LB1_line1, M4_CalP0_LP0_CL3_LB1_line2, M4_CalP0_LP0_CL3_line1);
or2 M4_CalP0_LP0_CL3_LB2(in389, M4_CalP0_LP0_CL3_line0, M4_CalP0_LP0_CL3_line2);
nand2 M4_CalP0_LP0_CL3_LB3(in389, M4_CalP0_LP0_CL3_line1, M4_CalP0_LP0_CL3_line3);
and2 M4_CalP0_LP0_CL3_LB4(M4_CalP0_LP0_CL3_line2, M4_CalP0_LP0_CL3_line3, M4_CalP0_LogicOut_3);
inv M4_CalP0_LP0_CL4_LB0_Mux2_0(in234, M4_CalP0_LP0_CL4_LB0_Not_ContIn);
and2 M4_CalP0_LP0_CL4_LB0_Mux2_1(in254, M4_CalP0_LP0_CL4_LB0_Not_ContIn, M4_CalP0_LP0_CL4_LB0_line1);
and2 M4_CalP0_LP0_CL4_LB0_Mux2_2(in242, in234, M4_CalP0_LP0_CL4_LB0_line2);
or2 M4_CalP0_LP0_CL4_LB0_Mux2_3(M4_CalP0_LP0_CL4_LB0_line1, M4_CalP0_LP0_CL4_LB0_line2, M4_CalP0_LP0_CL4_line0);
inv M4_CalP0_LP0_CL4_LB1_Mux2_0(in234, M4_CalP0_LP0_CL4_LB1_Not_ContIn);
and2 M4_CalP0_LP0_CL4_LB1_Mux2_1(in251, M4_CalP0_LP0_CL4_LB1_Not_ContIn, M4_CalP0_LP0_CL4_LB1_line1);
and2 M4_CalP0_LP0_CL4_LB1_Mux2_2(in248, in234, M4_CalP0_LP0_CL4_LB1_line2);
or2 M4_CalP0_LP0_CL4_LB1_Mux2_3(M4_CalP0_LP0_CL4_LB1_line1, M4_CalP0_LP0_CL4_LB1_line2, M4_CalP0_LP0_CL4_line1);
or2 M4_CalP0_LP0_CL4_LB2(in435, M4_CalP0_LP0_CL4_line0, M4_CalP0_LP0_CL4_line2);
nand2 M4_CalP0_LP0_CL4_LB3(in435, M4_CalP0_LP0_CL4_line1, M4_CalP0_LP0_CL4_line3);
and2 M4_CalP0_LP0_CL4_LB4(M4_CalP0_LP0_CL4_line2, M4_CalP0_LP0_CL4_line3, M4_CalP0_LogicOut_4);
inv M4_CalP0_LP0_CL5_LB0_Mux2_0(in226, M4_CalP0_LP0_CL5_LB0_Not_ContIn);
and2 M4_CalP0_LP0_CL5_LB0_Mux2_1(in254, M4_CalP0_LP0_CL5_LB0_Not_ContIn, M4_CalP0_LP0_CL5_LB0_line1);
and2 M4_CalP0_LP0_CL5_LB0_Mux2_2(in242, in226, M4_CalP0_LP0_CL5_LB0_line2);
or2 M4_CalP0_LP0_CL5_LB0_Mux2_3(M4_CalP0_LP0_CL5_LB0_line1, M4_CalP0_LP0_CL5_LB0_line2, M4_CalP0_LP0_CL5_line0);
inv M4_CalP0_LP0_CL5_LB1_Mux2_0(in226, M4_CalP0_LP0_CL5_LB1_Not_ContIn);
and2 M4_CalP0_LP0_CL5_LB1_Mux2_1(in251, M4_CalP0_LP0_CL5_LB1_Not_ContIn, M4_CalP0_LP0_CL5_LB1_line1);
and2 M4_CalP0_LP0_CL5_LB1_Mux2_2(in248, in226, M4_CalP0_LP0_CL5_LB1_line2);
or2 M4_CalP0_LP0_CL5_LB1_Mux2_3(M4_CalP0_LP0_CL5_LB1_line1, M4_CalP0_LP0_CL5_LB1_line2, M4_CalP0_LP0_CL5_line1);
or2 M4_CalP0_LP0_CL5_LB2(in422, M4_CalP0_LP0_CL5_line0, M4_CalP0_LP0_CL5_line2);
nand2 M4_CalP0_LP0_CL5_LB3(in422, M4_CalP0_LP0_CL5_line1, M4_CalP0_LP0_CL5_line3);
and2 M4_CalP0_LP0_CL5_LB4(M4_CalP0_LP0_CL5_line2, M4_CalP0_LP0_CL5_line3, M4_CalP0_LogicOut_5);
inv M4_CalP0_LP0_CL6_LB0_Mux2_0(in218, M4_CalP0_LP0_CL6_LB0_Not_ContIn);
and2 M4_CalP0_LP0_CL6_LB0_Mux2_1(in254, M4_CalP0_LP0_CL6_LB0_Not_ContIn, M4_CalP0_LP0_CL6_LB0_line1);
and2 M4_CalP0_LP0_CL6_LB0_Mux2_2(in242, in218, M4_CalP0_LP0_CL6_LB0_line2);
or2 M4_CalP0_LP0_CL6_LB0_Mux2_3(M4_CalP0_LP0_CL6_LB0_line1, M4_CalP0_LP0_CL6_LB0_line2, M4_CalP0_LP0_CL6_line0);
inv M4_CalP0_LP0_CL6_LB1_Mux2_0(in218, M4_CalP0_LP0_CL6_LB1_Not_ContIn);
and2 M4_CalP0_LP0_CL6_LB1_Mux2_1(in251, M4_CalP0_LP0_CL6_LB1_Not_ContIn, M4_CalP0_LP0_CL6_LB1_line1);
and2 M4_CalP0_LP0_CL6_LB1_Mux2_2(in248, in218, M4_CalP0_LP0_CL6_LB1_line2);
or2 M4_CalP0_LP0_CL6_LB1_Mux2_3(M4_CalP0_LP0_CL6_LB1_line1, M4_CalP0_LP0_CL6_LB1_line2, M4_CalP0_LP0_CL6_line1);
or2 M4_CalP0_LP0_CL6_LB2(in468, M4_CalP0_LP0_CL6_line0, M4_CalP0_LP0_CL6_line2);
nand2 M4_CalP0_LP0_CL6_LB3(in468, M4_CalP0_LP0_CL6_line1, M4_CalP0_LP0_CL6_line3);
and2 M4_CalP0_LP0_CL6_LB4(M4_CalP0_LP0_CL6_line2, M4_CalP0_LP0_CL6_line3, M4_CalP0_LogicOut_6);
inv M4_CalP0_LP0_CL7_LB0_Mux2_0(in210, M4_CalP0_LP0_CL7_LB0_Not_ContIn);
and2 M4_CalP0_LP0_CL7_LB0_Mux2_1(in254, M4_CalP0_LP0_CL7_LB0_Not_ContIn, M4_CalP0_LP0_CL7_LB0_line1);
and2 M4_CalP0_LP0_CL7_LB0_Mux2_2(in242, in210, M4_CalP0_LP0_CL7_LB0_line2);
or2 M4_CalP0_LP0_CL7_LB0_Mux2_3(M4_CalP0_LP0_CL7_LB0_line1, M4_CalP0_LP0_CL7_LB0_line2, M4_CalP0_LP0_CL7_line0);
inv M4_CalP0_LP0_CL7_LB1_Mux2_0(in210, M4_CalP0_LP0_CL7_LB1_Not_ContIn);
and2 M4_CalP0_LP0_CL7_LB1_Mux2_1(in251, M4_CalP0_LP0_CL7_LB1_Not_ContIn, M4_CalP0_LP0_CL7_LB1_line1);
and2 M4_CalP0_LP0_CL7_LB1_Mux2_2(in248, in210, M4_CalP0_LP0_CL7_LB1_line2);
or2 M4_CalP0_LP0_CL7_LB1_Mux2_3(M4_CalP0_LP0_CL7_LB1_line1, M4_CalP0_LP0_CL7_LB1_line2, M4_CalP0_LP0_CL7_line1);
or2 M4_CalP0_LP0_CL7_LB2(in457, M4_CalP0_LP0_CL7_line0, M4_CalP0_LP0_CL7_line2);
nand2 M4_CalP0_LP0_CL7_LB3(in457, M4_CalP0_LP0_CL7_line1, M4_CalP0_LP0_CL7_line3);
and2 M4_CalP0_LP0_CL7_LB4(M4_CalP0_LP0_CL7_line2, M4_CalP0_LP0_CL7_line3, M4_CalP0_LogicOut_7);
inv M4_CalP0_LP0_CL8_LB0_Mux2_0(in206, M4_CalP0_LP0_CL8_LB0_Not_ContIn);
and2 M4_CalP0_LP0_CL8_LB0_Mux2_1(in254, M4_CalP0_LP0_CL8_LB0_Not_ContIn, M4_CalP0_LP0_CL8_LB0_line1);
and2 M4_CalP0_LP0_CL8_LB0_Mux2_2(in242, in206, M4_CalP0_LP0_CL8_LB0_line2);
or2 M4_CalP0_LP0_CL8_LB0_Mux2_3(M4_CalP0_LP0_CL8_LB0_line1, M4_CalP0_LP0_CL8_LB0_line2, M4_CalP0_LP0_CL8_line0);
inv M4_CalP0_LP0_CL8_LB1_Mux2_0(in206, M4_CalP0_LP0_CL8_LB1_Not_ContIn);
and2 M4_CalP0_LP0_CL8_LB1_Mux2_1(in251, M4_CalP0_LP0_CL8_LB1_Not_ContIn, M4_CalP0_LP0_CL8_LB1_line1);
and2 M4_CalP0_LP0_CL8_LB1_Mux2_2(in248, in206, M4_CalP0_LP0_CL8_LB1_line2);
or2 M4_CalP0_LP0_CL8_LB1_Mux2_3(M4_CalP0_LP0_CL8_LB1_line1, M4_CalP0_LP0_CL8_LB1_line2, M4_CalP0_LP0_CL8_line1);
or2 M4_CalP0_LP0_CL8_LB2(in446, M4_CalP0_LP0_CL8_line0, M4_CalP0_LP0_CL8_line2);
nand2 M4_CalP0_LP0_CL8_LB3(in446, M4_CalP0_LP0_CL8_line1, M4_CalP0_LP0_CL8_line3);
and2 M4_CalP0_LP0_CL8_LB4(M4_CalP0_LP0_CL8_line2, M4_CalP0_LP0_CL8_line3, M4_CalP0_LogicOut_8);
inv M4_CalP0_LP1_PT1_Xo0(M4_CalP0_LogicOut_5, M4_CalP0_LP1_PT1_NotA);
inv M4_CalP0_LP1_PT1_Xo1(M4_CalP0_LogicOut_6, M4_CalP0_LP1_PT1_NotB);
nand2 M4_CalP0_LP1_PT1_Xo2(M4_CalP0_LP1_PT1_NotA, M4_CalP0_LogicOut_6, M4_CalP0_LP1_PT1_line2);
nand2 M4_CalP0_LP1_PT1_Xo3(M4_CalP0_LP1_PT1_NotB, M4_CalP0_LogicOut_5, M4_CalP0_LP1_PT1_line3);
nand2 M4_CalP0_LP1_PT1_Xo4(M4_CalP0_LP1_PT1_line2, M4_CalP0_LP1_PT1_line3, M4_CalP0_LP1_line1);
inv M4_CalP0_LP1_PT2_Xo0(M4_CalP0_LogicOut_7, M4_CalP0_LP1_PT2_NotA);
inv M4_CalP0_LP1_PT2_Xo1(M4_CalP0_LogicOut_8, M4_CalP0_LP1_PT2_NotB);
nand2 M4_CalP0_LP1_PT2_Xo2(M4_CalP0_LP1_PT2_NotA, M4_CalP0_LogicOut_8, M4_CalP0_LP1_PT2_line2);
nand2 M4_CalP0_LP1_PT2_Xo3(M4_CalP0_LP1_PT2_NotB, M4_CalP0_LogicOut_7, M4_CalP0_LP1_PT2_line3);
nand2 M4_CalP0_LP1_PT2_Xo4(M4_CalP0_LP1_PT2_line2, M4_CalP0_LP1_PT2_line3, M4_CalP0_LP1_line2);
inv M4_CalP0_LP1_PT3_Xo0(M4_CalP0_LogicOut_1, M4_CalP0_LP1_PT3_NotA);
inv M4_CalP0_LP1_PT3_Xo1(M4_CalP0_LogicOut_2, M4_CalP0_LP1_PT3_NotB);
nand2 M4_CalP0_LP1_PT3_Xo2(M4_CalP0_LP1_PT3_NotA, M4_CalP0_LogicOut_2, M4_CalP0_LP1_PT3_line2);
nand2 M4_CalP0_LP1_PT3_Xo3(M4_CalP0_LP1_PT3_NotB, M4_CalP0_LogicOut_1, M4_CalP0_LP1_PT3_line3);
nand2 M4_CalP0_LP1_PT3_Xo4(M4_CalP0_LP1_PT3_line2, M4_CalP0_LP1_PT3_line3, M4_CalP0_LP1_line3);
inv M4_CalP0_LP1_PT4_Xo0(M4_CalP0_LogicOut_3, M4_CalP0_LP1_PT4_NotA);
inv M4_CalP0_LP1_PT4_Xo1(M4_CalP0_LogicOut_4, M4_CalP0_LP1_PT4_NotB);
nand2 M4_CalP0_LP1_PT4_Xo2(M4_CalP0_LP1_PT4_NotA, M4_CalP0_LogicOut_4, M4_CalP0_LP1_PT4_line2);
nand2 M4_CalP0_LP1_PT4_Xo3(M4_CalP0_LP1_PT4_NotB, M4_CalP0_LogicOut_3, M4_CalP0_LP1_PT4_line3);
nand2 M4_CalP0_LP1_PT4_Xo4(M4_CalP0_LP1_PT4_line2, M4_CalP0_LP1_PT4_line3, M4_CalP0_LP1_line4);
inv M4_CalP0_LP1_PT5_Xo0(M4_CalP0_LP1_line1, M4_CalP0_LP1_PT5_NotA);
inv M4_CalP0_LP1_PT5_Xo1(M4_CalP0_LP1_line2, M4_CalP0_LP1_PT5_NotB);
nand2 M4_CalP0_LP1_PT5_Xo2(M4_CalP0_LP1_PT5_NotA, M4_CalP0_LP1_line2, M4_CalP0_LP1_PT5_line2);
nand2 M4_CalP0_LP1_PT5_Xo3(M4_CalP0_LP1_PT5_NotB, M4_CalP0_LP1_line1, M4_CalP0_LP1_PT5_line3);
nand2 M4_CalP0_LP1_PT5_Xo4(M4_CalP0_LP1_PT5_line2, M4_CalP0_LP1_PT5_line3, M4_CalP0_LP1_line5);
inv M4_CalP0_LP1_PT6_Xo3_0(M4_CalP0_LP1_line3, M4_CalP0_LP1_PT6_NotA);
inv M4_CalP0_LP1_PT6_Xo3_1(M4_CalP0_LogicOut_0, M4_CalP0_LP1_PT6_NotB);
inv M4_CalP0_LP1_PT6_Xo3_2(M4_CalP0_LP1_line4, M4_CalP0_LP1_PT6_NotC);
and3 M4_CalP0_LP1_PT6_Xo3_3(M4_CalP0_LP1_PT6_NotA, M4_CalP0_LP1_PT6_NotB, M4_CalP0_LP1_line4, M4_CalP0_LP1_PT6_line3);
and3 M4_CalP0_LP1_PT6_Xo3_4(M4_CalP0_LP1_PT6_NotA, M4_CalP0_LogicOut_0, M4_CalP0_LP1_PT6_NotC, M4_CalP0_LP1_PT6_line4);
and3 M4_CalP0_LP1_PT6_Xo3_5(M4_CalP0_LP1_line3, M4_CalP0_LP1_PT6_NotB, M4_CalP0_LP1_PT6_NotC, M4_CalP0_LP1_PT6_line5);
and3 M4_CalP0_LP1_PT6_Xo3_6(M4_CalP0_LP1_line3, M4_CalP0_LogicOut_0, M4_CalP0_LP1_line4, M4_CalP0_LP1_PT6_line6);
nor2 M4_CalP0_LP1_PT6_Xo3_7(M4_CalP0_LP1_PT6_line3, M4_CalP0_LP1_PT6_line4, M4_CalP0_LP1_PT6_line7);
nor2 M4_CalP0_LP1_PT6_Xo3_8(M4_CalP0_LP1_PT6_line5, M4_CalP0_LP1_PT6_line6, M4_CalP0_LP1_PT6_line8);
nand2 M4_CalP0_LP1_PT6_Xo3_9(M4_CalP0_LP1_PT6_line7, M4_CalP0_LP1_PT6_line8, M4_CalP0_LP1_line6);
inv M4_CalP0_LP1_PT7_Xo0(M4_CalP0_LP1_line5, M4_CalP0_LP1_PT7_NotA);
inv M4_CalP0_LP1_PT7_Xo1(M4_CalP0_LP1_line6, M4_CalP0_LP1_PT7_NotB);
nand2 M4_CalP0_LP1_PT7_Xo2(M4_CalP0_LP1_PT7_NotA, M4_CalP0_LP1_line6, M4_CalP0_LP1_PT7_line2);
nand2 M4_CalP0_LP1_PT7_Xo3(M4_CalP0_LP1_PT7_NotB, M4_CalP0_LP1_line5, M4_CalP0_LP1_PT7_line3);
nand2 M4_CalP0_LP1_PT7_Xo4(M4_CalP0_LP1_PT7_line2, M4_CalP0_LP1_PT7_line3, M4_LogicPar);
and2 M4_CalP1_SP0_GP9_0(Ybus_0, in374, M4_CalP1_Genbus_0);
and2 M4_CalP1_SP0_GP9_1(Ybus_1, in411, M4_CalP1_Genbus_1);
and2 M4_CalP1_SP0_GP9_2(Ybus_2, in400, M4_CalP1_Genbus_2);
and2 M4_CalP1_SP0_GP9_3(Ybus_3, in389, M4_CalP1_Genbus_3);
and2 M4_CalP1_SP0_GP9_4(Ybus_4, in435, M4_CalP1_Genbus_4);
and2 M4_CalP1_SP0_GP9_5(Ybus_5, in422, M4_CalP1_Genbus_5);
and2 M4_CalP1_SP0_GP9_6(Ybus_6, in468, M4_CalP1_Genbus_6);
and2 M4_CalP1_SP0_GP9_7(Ybus_7, in457, M4_CalP1_Genbus_7);
and2 M4_CalP1_SP0_GP9_8(Ybus_8, in446, M4_CalP1_Genbus_8);
inv M4_CalP1_SP0_GP9_9_Xo0(Ybus_0, M4_CalP1_SP0_GP9_9_NotA);
inv M4_CalP1_SP0_GP9_9_Xo1(in374, M4_CalP1_SP0_GP9_9_NotB);
nand2 M4_CalP1_SP0_GP9_9_Xo2(M4_CalP1_SP0_GP9_9_NotA, in374, M4_CalP1_SP0_GP9_9_line2);
nand2 M4_CalP1_SP0_GP9_9_Xo3(M4_CalP1_SP0_GP9_9_NotB, Ybus_0, M4_CalP1_SP0_GP9_9_line3);
nand2 M4_CalP1_SP0_GP9_9_Xo4(M4_CalP1_SP0_GP9_9_line2, M4_CalP1_SP0_GP9_9_line3, M4_CalP1_Propbus_0);
inv M4_CalP1_SP0_GP9_10_Xo0(Ybus_1, M4_CalP1_SP0_GP9_10_NotA);
inv M4_CalP1_SP0_GP9_10_Xo1(in411, M4_CalP1_SP0_GP9_10_NotB);
nand2 M4_CalP1_SP0_GP9_10_Xo2(M4_CalP1_SP0_GP9_10_NotA, in411, M4_CalP1_SP0_GP9_10_line2);
nand2 M4_CalP1_SP0_GP9_10_Xo3(M4_CalP1_SP0_GP9_10_NotB, Ybus_1, M4_CalP1_SP0_GP9_10_line3);
nand2 M4_CalP1_SP0_GP9_10_Xo4(M4_CalP1_SP0_GP9_10_line2, M4_CalP1_SP0_GP9_10_line3, M4_CalP1_Propbus_1);
inv M4_CalP1_SP0_GP9_11_Xo0(Ybus_2, M4_CalP1_SP0_GP9_11_NotA);
inv M4_CalP1_SP0_GP9_11_Xo1(in400, M4_CalP1_SP0_GP9_11_NotB);
nand2 M4_CalP1_SP0_GP9_11_Xo2(M4_CalP1_SP0_GP9_11_NotA, in400, M4_CalP1_SP0_GP9_11_line2);
nand2 M4_CalP1_SP0_GP9_11_Xo3(M4_CalP1_SP0_GP9_11_NotB, Ybus_2, M4_CalP1_SP0_GP9_11_line3);
nand2 M4_CalP1_SP0_GP9_11_Xo4(M4_CalP1_SP0_GP9_11_line2, M4_CalP1_SP0_GP9_11_line3, M4_CalP1_Propbus_2);
inv M4_CalP1_SP0_GP9_12_Xo0(Ybus_3, M4_CalP1_SP0_GP9_12_NotA);
inv M4_CalP1_SP0_GP9_12_Xo1(in389, M4_CalP1_SP0_GP9_12_NotB);
nand2 M4_CalP1_SP0_GP9_12_Xo2(M4_CalP1_SP0_GP9_12_NotA, in389, M4_CalP1_SP0_GP9_12_line2);
nand2 M4_CalP1_SP0_GP9_12_Xo3(M4_CalP1_SP0_GP9_12_NotB, Ybus_3, M4_CalP1_SP0_GP9_12_line3);
nand2 M4_CalP1_SP0_GP9_12_Xo4(M4_CalP1_SP0_GP9_12_line2, M4_CalP1_SP0_GP9_12_line3, M4_CalP1_Propbus_3);
inv M4_CalP1_SP0_GP9_13_Xo0(Ybus_4, M4_CalP1_SP0_GP9_13_NotA);
inv M4_CalP1_SP0_GP9_13_Xo1(in435, M4_CalP1_SP0_GP9_13_NotB);
nand2 M4_CalP1_SP0_GP9_13_Xo2(M4_CalP1_SP0_GP9_13_NotA, in435, M4_CalP1_SP0_GP9_13_line2);
nand2 M4_CalP1_SP0_GP9_13_Xo3(M4_CalP1_SP0_GP9_13_NotB, Ybus_4, M4_CalP1_SP0_GP9_13_line3);
nand2 M4_CalP1_SP0_GP9_13_Xo4(M4_CalP1_SP0_GP9_13_line2, M4_CalP1_SP0_GP9_13_line3, M4_CalP1_Propbus_4);
inv M4_CalP1_SP0_GP9_14_Xo0(Ybus_5, M4_CalP1_SP0_GP9_14_NotA);
inv M4_CalP1_SP0_GP9_14_Xo1(in422, M4_CalP1_SP0_GP9_14_NotB);
nand2 M4_CalP1_SP0_GP9_14_Xo2(M4_CalP1_SP0_GP9_14_NotA, in422, M4_CalP1_SP0_GP9_14_line2);
nand2 M4_CalP1_SP0_GP9_14_Xo3(M4_CalP1_SP0_GP9_14_NotB, Ybus_5, M4_CalP1_SP0_GP9_14_line3);
nand2 M4_CalP1_SP0_GP9_14_Xo4(M4_CalP1_SP0_GP9_14_line2, M4_CalP1_SP0_GP9_14_line3, M4_CalP1_Propbus_5);
inv M4_CalP1_SP0_GP9_15_Xo0(Ybus_6, M4_CalP1_SP0_GP9_15_NotA);
inv M4_CalP1_SP0_GP9_15_Xo1(in468, M4_CalP1_SP0_GP9_15_NotB);
nand2 M4_CalP1_SP0_GP9_15_Xo2(M4_CalP1_SP0_GP9_15_NotA, in468, M4_CalP1_SP0_GP9_15_line2);
nand2 M4_CalP1_SP0_GP9_15_Xo3(M4_CalP1_SP0_GP9_15_NotB, Ybus_6, M4_CalP1_SP0_GP9_15_line3);
nand2 M4_CalP1_SP0_GP9_15_Xo4(M4_CalP1_SP0_GP9_15_line2, M4_CalP1_SP0_GP9_15_line3, M4_CalP1_Propbus_6);
inv M4_CalP1_SP0_GP9_16_Xo0(Ybus_7, M4_CalP1_SP0_GP9_16_NotA);
inv M4_CalP1_SP0_GP9_16_Xo1(in457, M4_CalP1_SP0_GP9_16_NotB);
nand2 M4_CalP1_SP0_GP9_16_Xo2(M4_CalP1_SP0_GP9_16_NotA, in457, M4_CalP1_SP0_GP9_16_line2);
nand2 M4_CalP1_SP0_GP9_16_Xo3(M4_CalP1_SP0_GP9_16_NotB, Ybus_7, M4_CalP1_SP0_GP9_16_line3);
nand2 M4_CalP1_SP0_GP9_16_Xo4(M4_CalP1_SP0_GP9_16_line2, M4_CalP1_SP0_GP9_16_line3, M4_CalP1_Propbus_7);
inv M4_CalP1_SP0_GP9_17_Xo0(Ybus_8, M4_CalP1_SP0_GP9_17_NotA);
inv M4_CalP1_SP0_GP9_17_Xo1(in446, M4_CalP1_SP0_GP9_17_NotB);
nand2 M4_CalP1_SP0_GP9_17_Xo2(M4_CalP1_SP0_GP9_17_NotA, in446, M4_CalP1_SP0_GP9_17_line2);
nand2 M4_CalP1_SP0_GP9_17_Xo3(M4_CalP1_SP0_GP9_17_NotB, Ybus_8, M4_CalP1_SP0_GP9_17_line3);
nand2 M4_CalP1_SP0_GP9_17_Xo4(M4_CalP1_SP0_GP9_17_line2, M4_CalP1_SP0_GP9_17_line3, M4_CalP1_Propbus_8);
or2 M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_0(M4_CalP1_Genbus_0, M4_CalP1_Propbus_0, M4_CalP1_LocalC1_0);
and2 M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_1_Ao2_0(M4_CalP1_Propbus_1, M4_CalP1_Genbus_0, M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_1_line0);
or2 M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_1_Ao2_1(M4_CalP1_Genbus_1, M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_1_line0, M4_CalP1_LocalC0_1);
and2 M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_2_Ao3a_0(M4_CalP1_Propbus_1, M4_CalP1_Genbus_0, M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_2_line0);
and2 M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_2_Ao3a_1(M4_CalP1_Propbus_1, M4_CalP1_Propbus_0, M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_2_line1);
or3 M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_2_Ao3a_2(M4_CalP1_Genbus_1, M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_2_line0, M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_2_line1, M4_CalP1_LocalC1_1);
and2 M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_3_Ao3a_0(M4_CalP1_Propbus_2, M4_CalP1_Genbus_1, M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_3_line0);
and3 M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_3_Ao3a_1(M4_CalP1_Propbus_2, M4_CalP1_Propbus_1, M4_CalP1_Genbus_0, M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_3_line1);
or3 M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_3_Ao3a_2(M4_CalP1_Genbus_2, M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_3_line0, M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_3_line1, M4_CalP1_LocalC0_2);
and2 M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_4_Ao4a_0(M4_CalP1_Propbus_2, M4_CalP1_Genbus_1, M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_4_line0);
and3 M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_4_Ao4a_1(M4_CalP1_Propbus_2, M4_CalP1_Propbus_1, M4_CalP1_Genbus_0, M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_4_line1);
and3 M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_4_Ao4a_2(M4_CalP1_Propbus_2, M4_CalP1_Propbus_1, M4_CalP1_Propbus_0, M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_4_line2);
or4 M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_4_Ao4a_3(M4_CalP1_Genbus_2, M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_4_line0, M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_4_line1, M4_CalP1_SP1_GLC5_0_GLC4_0_GLC4_4_line2, M4_CalP1_LocalC1_2);
and2 M4_CalP1_SP1_GLC5_0_GLC4_1_Ao4a_0(M4_CalP1_Propbus_3, M4_CalP1_Genbus_2, M4_CalP1_SP1_GLC5_0_GLC4_1_line0);
and3 M4_CalP1_SP1_GLC5_0_GLC4_1_Ao4a_1(M4_CalP1_Propbus_3, M4_CalP1_Propbus_2, M4_CalP1_Genbus_1, M4_CalP1_SP1_GLC5_0_GLC4_1_line1);
and4 M4_CalP1_SP1_GLC5_0_GLC4_1_Ao4a_2(M4_CalP1_Propbus_3, M4_CalP1_Propbus_2, M4_CalP1_Propbus_1, M4_CalP1_Genbus_0, M4_CalP1_SP1_GLC5_0_GLC4_1_line2);
or4 M4_CalP1_SP1_GLC5_0_GLC4_1_Ao4a_3(M4_CalP1_Genbus_3, M4_CalP1_SP1_GLC5_0_GLC4_1_line0, M4_CalP1_SP1_GLC5_0_GLC4_1_line1, M4_CalP1_SP1_GLC5_0_GLC4_1_line2, M4_CalP1_LocalC0_3);
and2 M4_CalP1_SP1_GLC5_0_GLC4_2_Ao5a_0(M4_CalP1_Propbus_3, M4_CalP1_Genbus_2, M4_CalP1_SP1_GLC5_0_GLC4_2_line0);
and3 M4_CalP1_SP1_GLC5_0_GLC4_2_Ao5a_1(M4_CalP1_Propbus_3, M4_CalP1_Propbus_2, M4_CalP1_Genbus_1, M4_CalP1_SP1_GLC5_0_GLC4_2_line1);
and4 M4_CalP1_SP1_GLC5_0_GLC4_2_Ao5a_2(M4_CalP1_Propbus_3, M4_CalP1_Propbus_2, M4_CalP1_Propbus_1, M4_CalP1_Genbus_0, M4_CalP1_SP1_GLC5_0_GLC4_2_line2);
and4 M4_CalP1_SP1_GLC5_0_GLC4_2_Ao5a_3(M4_CalP1_Propbus_3, M4_CalP1_Propbus_2, M4_CalP1_Propbus_1, M4_CalP1_Propbus_0, M4_CalP1_SP1_GLC5_0_GLC4_2_line3);
or5 M4_CalP1_SP1_GLC5_0_GLC4_2_Ao5a_4(M4_CalP1_Genbus_3, M4_CalP1_SP1_GLC5_0_GLC4_2_line0, M4_CalP1_SP1_GLC5_0_GLC4_2_line1, M4_CalP1_SP1_GLC5_0_GLC4_2_line2, M4_CalP1_SP1_GLC5_0_GLC4_2_line3, M4_CalP1_LocalC1_3);
and2 M4_CalP1_SP1_GLC5_1_Ao5a_0(M4_CalP1_Propbus_4, M4_CalP1_Genbus_3, M4_CalP1_SP1_GLC5_1_line0);
and3 M4_CalP1_SP1_GLC5_1_Ao5a_1(M4_CalP1_Propbus_4, M4_CalP1_Propbus_3, M4_CalP1_Genbus_2, M4_CalP1_SP1_GLC5_1_line1);
and4 M4_CalP1_SP1_GLC5_1_Ao5a_2(M4_CalP1_Propbus_4, M4_CalP1_Propbus_3, M4_CalP1_Propbus_2, M4_CalP1_Genbus_1, M4_CalP1_SP1_GLC5_1_line2);
and5 M4_CalP1_SP1_GLC5_1_Ao5a_3(M4_CalP1_Propbus_4, M4_CalP1_Propbus_3, M4_CalP1_Propbus_2, M4_CalP1_Propbus_1, M4_CalP1_Genbus_0, M4_CalP1_SP1_GLC5_1_line3);
or5 M4_CalP1_SP1_GLC5_1_Ao5a_4(M4_CalP1_Genbus_4, M4_CalP1_SP1_GLC5_1_line0, M4_CalP1_SP1_GLC5_1_line1, M4_CalP1_SP1_GLC5_1_line2, M4_CalP1_SP1_GLC5_1_line3, M4_CalP1_LocalC0_4);
and2 M4_CalP1_SP1_GLC5_2_Ao6a_0(M4_CalP1_Propbus_4, M4_CalP1_Genbus_3, M4_CalP1_SP1_GLC5_2_line0);
and3 M4_CalP1_SP1_GLC5_2_Ao6a_1(M4_CalP1_Propbus_4, M4_CalP1_Propbus_3, M4_CalP1_Genbus_2, M4_CalP1_SP1_GLC5_2_line1);
and4 M4_CalP1_SP1_GLC5_2_Ao6a_2(M4_CalP1_Propbus_4, M4_CalP1_Propbus_3, M4_CalP1_Propbus_2, M4_CalP1_Genbus_1, M4_CalP1_SP1_GLC5_2_line2);
and5 M4_CalP1_SP1_GLC5_2_Ao6a_3(M4_CalP1_Propbus_4, M4_CalP1_Propbus_3, M4_CalP1_Propbus_2, M4_CalP1_Propbus_1, M4_CalP1_Genbus_0, M4_CalP1_SP1_GLC5_2_line3);
and5 M4_CalP1_SP1_GLC5_2_Ao6a_4(M4_CalP1_Propbus_4, M4_CalP1_Propbus_3, M4_CalP1_Propbus_2, M4_CalP1_Propbus_1, M4_CalP1_Propbus_0, M4_CalP1_SP1_GLC5_2_line4);
or6 M4_CalP1_SP1_GLC5_2_Ao6a_5(M4_CalP1_Genbus_4, M4_CalP1_SP1_GLC5_2_line0, M4_CalP1_SP1_GLC5_2_line1, M4_CalP1_SP1_GLC5_2_line2, M4_CalP1_SP1_GLC5_2_line3, M4_CalP1_SP1_GLC5_2_line4, M4_CalP1_LocalC1_4);
or2 M4_CalP1_SP2_GLC4_0(M4_CalP1_Genbus_5, M4_CalP1_Propbus_5, M4_CalP1_LocalC1_5);
and2 M4_CalP1_SP2_GLC4_1_Ao2_0(M4_CalP1_Propbus_6, M4_CalP1_Genbus_5, M4_CalP1_SP2_GLC4_1_line0);
or2 M4_CalP1_SP2_GLC4_1_Ao2_1(M4_CalP1_Genbus_6, M4_CalP1_SP2_GLC4_1_line0, M4_CalP1_LocalC0_6);
and2 M4_CalP1_SP2_GLC4_2_Ao3a_0(M4_CalP1_Propbus_6, M4_CalP1_Genbus_5, M4_CalP1_SP2_GLC4_2_line0);
and2 M4_CalP1_SP2_GLC4_2_Ao3a_1(M4_CalP1_Propbus_6, M4_CalP1_Propbus_5, M4_CalP1_SP2_GLC4_2_line1);
or3 M4_CalP1_SP2_GLC4_2_Ao3a_2(M4_CalP1_Genbus_6, M4_CalP1_SP2_GLC4_2_line0, M4_CalP1_SP2_GLC4_2_line1, M4_CalP1_LocalC1_6);
and2 M4_CalP1_SP2_GLC4_3_Ao3a_0(M4_CalP1_Propbus_7, M4_CalP1_Genbus_6, M4_CalP1_SP2_GLC4_3_line0);
and3 M4_CalP1_SP2_GLC4_3_Ao3a_1(M4_CalP1_Propbus_7, M4_CalP1_Propbus_6, M4_CalP1_Genbus_5, M4_CalP1_SP2_GLC4_3_line1);
or3 M4_CalP1_SP2_GLC4_3_Ao3a_2(M4_CalP1_Genbus_7, M4_CalP1_SP2_GLC4_3_line0, M4_CalP1_SP2_GLC4_3_line1, M4_CalP1_LocalC0_7);
and2 M4_CalP1_SP2_GLC4_4_Ao4a_0(M4_CalP1_Propbus_7, M4_CalP1_Genbus_6, M4_CalP1_SP2_GLC4_4_line0);
and3 M4_CalP1_SP2_GLC4_4_Ao4a_1(M4_CalP1_Propbus_7, M4_CalP1_Propbus_6, M4_CalP1_Genbus_5, M4_CalP1_SP2_GLC4_4_line1);
and3 M4_CalP1_SP2_GLC4_4_Ao4a_2(M4_CalP1_Propbus_7, M4_CalP1_Propbus_6, M4_CalP1_Propbus_5, M4_CalP1_SP2_GLC4_4_line2);
or4 M4_CalP1_SP2_GLC4_4_Ao4a_3(M4_CalP1_Genbus_7, M4_CalP1_SP2_GLC4_4_line0, M4_CalP1_SP2_GLC4_4_line1, M4_CalP1_SP2_GLC4_4_line2, M4_CalP1_LocalC1_7);
inv M4_CalP1_SP3_SP9nc0_SP7nc0_Xo0(M4_CalP1_Genbus_0, M4_CalP1_SP3_SP9nc0_SP7nc0_NotA);
inv M4_CalP1_SP3_SP9nc0_SP7nc0_Xo1(M4_CalP1_LocalC0_1, M4_CalP1_SP3_SP9nc0_SP7nc0_NotB);
nand2 M4_CalP1_SP3_SP9nc0_SP7nc0_Xo2(M4_CalP1_SP3_SP9nc0_SP7nc0_NotA, M4_CalP1_LocalC0_1, M4_CalP1_SP3_SP9nc0_SP7nc0_line2);
nand2 M4_CalP1_SP3_SP9nc0_SP7nc0_Xo3(M4_CalP1_SP3_SP9nc0_SP7nc0_NotB, M4_CalP1_Genbus_0, M4_CalP1_SP3_SP9nc0_SP7nc0_line3);
nand2 M4_CalP1_SP3_SP9nc0_SP7nc0_Xo4(M4_CalP1_SP3_SP9nc0_SP7nc0_line2, M4_CalP1_SP3_SP9nc0_SP7nc0_line3, M4_CalP1_SP3_SP9nc0_line0);
inv M4_CalP1_SP3_SP9nc0_SP7nc1_Xo0(M4_CalP1_LocalC0_2, M4_CalP1_SP3_SP9nc0_SP7nc1_NotA);
inv M4_CalP1_SP3_SP9nc0_SP7nc1_Xo1(M4_CalP1_SP3_SP9nc0_line0, M4_CalP1_SP3_SP9nc0_SP7nc1_NotB);
nand2 M4_CalP1_SP3_SP9nc0_SP7nc1_Xo2(M4_CalP1_SP3_SP9nc0_SP7nc1_NotA, M4_CalP1_SP3_SP9nc0_line0, M4_CalP1_SP3_SP9nc0_SP7nc1_line2);
nand2 M4_CalP1_SP3_SP9nc0_SP7nc1_Xo3(M4_CalP1_SP3_SP9nc0_SP7nc1_NotB, M4_CalP1_LocalC0_2, M4_CalP1_SP3_SP9nc0_SP7nc1_line3);
nand2 M4_CalP1_SP3_SP9nc0_SP7nc1_Xo4(M4_CalP1_SP3_SP9nc0_SP7nc1_line2, M4_CalP1_SP3_SP9nc0_SP7nc1_line3, M4_CalP1_SP3_SP9nc0_line1);
inv M4_CalP1_SP3_SP9nc0_SP7nc2_Xo0(M4_CalP1_LocalC0_3, M4_CalP1_SP3_SP9nc0_SP7nc2_NotA);
inv M4_CalP1_SP3_SP9nc0_SP7nc2_Xo1(M4_CalP1_SP3_SP9nc0_line1, M4_CalP1_SP3_SP9nc0_SP7nc2_NotB);
nand2 M4_CalP1_SP3_SP9nc0_SP7nc2_Xo2(M4_CalP1_SP3_SP9nc0_SP7nc2_NotA, M4_CalP1_SP3_SP9nc0_line1, M4_CalP1_SP3_SP9nc0_SP7nc2_line2);
nand2 M4_CalP1_SP3_SP9nc0_SP7nc2_Xo3(M4_CalP1_SP3_SP9nc0_SP7nc2_NotB, M4_CalP1_LocalC0_3, M4_CalP1_SP3_SP9nc0_SP7nc2_line3);
nand2 M4_CalP1_SP3_SP9nc0_SP7nc2_Xo4(M4_CalP1_SP3_SP9nc0_SP7nc2_line2, M4_CalP1_SP3_SP9nc0_SP7nc2_line3, M4_CalP1_SP3_SP9nc0_line2);
inv M4_CalP1_SP3_SP9nc0_SP7nc3_Xo0(M4_CalP1_Propbus_0, M4_CalP1_SP3_SP9nc0_SP7nc3_NotA);
inv M4_CalP1_SP3_SP9nc0_SP7nc3_Xo1(M4_CalP1_SP3_SP9nc0_line2, M4_CalP1_SP3_SP9nc0_SP7nc3_NotB);
nand2 M4_CalP1_SP3_SP9nc0_SP7nc3_Xo2(M4_CalP1_SP3_SP9nc0_SP7nc3_NotA, M4_CalP1_SP3_SP9nc0_line2, M4_CalP1_SP3_SP9nc0_SP7nc3_line2);
nand2 M4_CalP1_SP3_SP9nc0_SP7nc3_Xo3(M4_CalP1_SP3_SP9nc0_SP7nc3_NotB, M4_CalP1_Propbus_0, M4_CalP1_SP3_SP9nc0_SP7nc3_line3);
nand2 M4_CalP1_SP3_SP9nc0_SP7nc3_Xo4(M4_CalP1_SP3_SP9nc0_SP7nc3_line2, M4_CalP1_SP3_SP9nc0_SP7nc3_line3, M4_CalP1_SP3_SP9nc0_line3);
inv M4_CalP1_SP3_SP9nc0_SP7nc4_Xo0(M4_CalP1_Propbus_1, M4_CalP1_SP3_SP9nc0_SP7nc4_NotA);
inv M4_CalP1_SP3_SP9nc0_SP7nc4_Xo1(M4_CalP1_SP3_SP9nc0_line3, M4_CalP1_SP3_SP9nc0_SP7nc4_NotB);
nand2 M4_CalP1_SP3_SP9nc0_SP7nc4_Xo2(M4_CalP1_SP3_SP9nc0_SP7nc4_NotA, M4_CalP1_SP3_SP9nc0_line3, M4_CalP1_SP3_SP9nc0_SP7nc4_line2);
nand2 M4_CalP1_SP3_SP9nc0_SP7nc4_Xo3(M4_CalP1_SP3_SP9nc0_SP7nc4_NotB, M4_CalP1_Propbus_1, M4_CalP1_SP3_SP9nc0_SP7nc4_line3);
nand2 M4_CalP1_SP3_SP9nc0_SP7nc4_Xo4(M4_CalP1_SP3_SP9nc0_SP7nc4_line2, M4_CalP1_SP3_SP9nc0_SP7nc4_line3, M4_CalP1_SP3_SP9nc0_line4);
inv M4_CalP1_SP3_SP9nc0_SP7nc5_Xo0(M4_CalP1_Propbus_2, M4_CalP1_SP3_SP9nc0_SP7nc5_NotA);
inv M4_CalP1_SP3_SP9nc0_SP7nc5_Xo1(M4_CalP1_SP3_SP9nc0_line4, M4_CalP1_SP3_SP9nc0_SP7nc5_NotB);
nand2 M4_CalP1_SP3_SP9nc0_SP7nc5_Xo2(M4_CalP1_SP3_SP9nc0_SP7nc5_NotA, M4_CalP1_SP3_SP9nc0_line4, M4_CalP1_SP3_SP9nc0_SP7nc5_line2);
nand2 M4_CalP1_SP3_SP9nc0_SP7nc5_Xo3(M4_CalP1_SP3_SP9nc0_SP7nc5_NotB, M4_CalP1_Propbus_2, M4_CalP1_SP3_SP9nc0_SP7nc5_line3);
nand2 M4_CalP1_SP3_SP9nc0_SP7nc5_Xo4(M4_CalP1_SP3_SP9nc0_SP7nc5_line2, M4_CalP1_SP3_SP9nc0_SP7nc5_line3, M4_CalP1_SP3_line0);
inv M4_CalP1_SP3_SP9nc1_Xo0(M4_CalP1_Propbus_3, M4_CalP1_SP3_SP9nc1_NotA);
inv M4_CalP1_SP3_SP9nc1_Xo1(M4_CalP1_SP3_line0, M4_CalP1_SP3_SP9nc1_NotB);
nand2 M4_CalP1_SP3_SP9nc1_Xo2(M4_CalP1_SP3_SP9nc1_NotA, M4_CalP1_SP3_line0, M4_CalP1_SP3_SP9nc1_line2);
nand2 M4_CalP1_SP3_SP9nc1_Xo3(M4_CalP1_SP3_SP9nc1_NotB, M4_CalP1_Propbus_3, M4_CalP1_SP3_SP9nc1_line3);
nand2 M4_CalP1_SP3_SP9nc1_Xo4(M4_CalP1_SP3_SP9nc1_line2, M4_CalP1_SP3_SP9nc1_line3, M4_CalP1_SP3_line1);
inv M4_CalP1_SP3_SP9nc2_Xo0(M4_CalP1_Propbus_4, M4_CalP1_SP3_SP9nc2_NotA);
inv M4_CalP1_SP3_SP9nc2_Xo1(M4_CalP1_SP3_line1, M4_CalP1_SP3_SP9nc2_NotB);
nand2 M4_CalP1_SP3_SP9nc2_Xo2(M4_CalP1_SP3_SP9nc2_NotA, M4_CalP1_SP3_line1, M4_CalP1_SP3_SP9nc2_line2);
nand2 M4_CalP1_SP3_SP9nc2_Xo3(M4_CalP1_SP3_SP9nc2_NotB, M4_CalP1_Propbus_4, M4_CalP1_SP3_SP9nc2_line3);
nand2 M4_CalP1_SP3_SP9nc2_Xo4(M4_CalP1_SP3_SP9nc2_line2, M4_CalP1_SP3_SP9nc2_line3, M4_CalP1_ParLo0);
inv M4_CalP1_SP4_SP9nc0_SP7c0(M4_CalP1_Propbus_2, M4_CalP1_SP4_SP9nc0_NewInbus_6);
inv M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_Xo0(M4_CalP1_LocalC1_0, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_NotA);
inv M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_Xo1(M4_CalP1_LocalC1_1, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_NotB);
nand2 M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_Xo2(M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_NotA, M4_CalP1_LocalC1_1, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_line2);
nand2 M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_Xo3(M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_NotB, M4_CalP1_LocalC1_0, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_line3);
nand2 M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_Xo4(M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_line2, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc0_line3, M4_CalP1_SP4_SP9nc0_SP7c2_line0);
inv M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_Xo0(M4_CalP1_LocalC1_2, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_NotA);
inv M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_Xo1(M4_CalP1_SP4_SP9nc0_SP7c2_line0, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_NotB);
nand2 M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_Xo2(M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_NotA, M4_CalP1_SP4_SP9nc0_SP7c2_line0, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_line2);
nand2 M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_Xo3(M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_NotB, M4_CalP1_LocalC1_2, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_line3);
nand2 M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_Xo4(M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_line2, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc1_line3, M4_CalP1_SP4_SP9nc0_SP7c2_line1);
inv M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_Xo0(M4_CalP1_LocalC1_3, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_NotA);
inv M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_Xo1(M4_CalP1_SP4_SP9nc0_SP7c2_line1, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_NotB);
nand2 M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_Xo2(M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_NotA, M4_CalP1_SP4_SP9nc0_SP7c2_line1, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_line2);
nand2 M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_Xo3(M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_NotB, M4_CalP1_LocalC1_3, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_line3);
nand2 M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_Xo4(M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_line2, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc2_line3, M4_CalP1_SP4_SP9nc0_SP7c2_line2);
inv M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_Xo0(M4_CalP1_Propbus_0, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_NotA);
inv M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_Xo1(M4_CalP1_SP4_SP9nc0_SP7c2_line2, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_NotB);
nand2 M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_Xo2(M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_NotA, M4_CalP1_SP4_SP9nc0_SP7c2_line2, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_line2);
nand2 M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_Xo3(M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_NotB, M4_CalP1_Propbus_0, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_line3);
nand2 M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_Xo4(M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_line2, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc3_line3, M4_CalP1_SP4_SP9nc0_SP7c2_line3);
inv M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_Xo0(M4_CalP1_Propbus_1, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_NotA);
inv M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_Xo1(M4_CalP1_SP4_SP9nc0_SP7c2_line3, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_NotB);
nand2 M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_Xo2(M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_NotA, M4_CalP1_SP4_SP9nc0_SP7c2_line3, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_line2);
nand2 M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_Xo3(M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_NotB, M4_CalP1_Propbus_1, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_line3);
nand2 M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_Xo4(M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_line2, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc4_line3, M4_CalP1_SP4_SP9nc0_SP7c2_line4);
inv M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_Xo0(M4_CalP1_SP4_SP9nc0_NewInbus_6, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_NotA);
inv M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_Xo1(M4_CalP1_SP4_SP9nc0_SP7c2_line4, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_NotB);
nand2 M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_Xo2(M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_NotA, M4_CalP1_SP4_SP9nc0_SP7c2_line4, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_line2);
nand2 M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_Xo3(M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_NotB, M4_CalP1_SP4_SP9nc0_NewInbus_6, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_line3);
nand2 M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_Xo4(M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_line2, M4_CalP1_SP4_SP9nc0_SP7c2_SP7nc5_line3, M4_CalP1_SP4_line0);
inv M4_CalP1_SP4_SP9nc1_Xo0(M4_CalP1_Propbus_3, M4_CalP1_SP4_SP9nc1_NotA);
inv M4_CalP1_SP4_SP9nc1_Xo1(M4_CalP1_SP4_line0, M4_CalP1_SP4_SP9nc1_NotB);
nand2 M4_CalP1_SP4_SP9nc1_Xo2(M4_CalP1_SP4_SP9nc1_NotA, M4_CalP1_SP4_line0, M4_CalP1_SP4_SP9nc1_line2);
nand2 M4_CalP1_SP4_SP9nc1_Xo3(M4_CalP1_SP4_SP9nc1_NotB, M4_CalP1_Propbus_3, M4_CalP1_SP4_SP9nc1_line3);
nand2 M4_CalP1_SP4_SP9nc1_Xo4(M4_CalP1_SP4_SP9nc1_line2, M4_CalP1_SP4_SP9nc1_line3, M4_CalP1_SP4_line1);
inv M4_CalP1_SP4_SP9nc2_Xo0(M4_CalP1_Propbus_4, M4_CalP1_SP4_SP9nc2_NotA);
inv M4_CalP1_SP4_SP9nc2_Xo1(M4_CalP1_SP4_line1, M4_CalP1_SP4_SP9nc2_NotB);
nand2 M4_CalP1_SP4_SP9nc2_Xo2(M4_CalP1_SP4_SP9nc2_NotA, M4_CalP1_SP4_line1, M4_CalP1_SP4_SP9nc2_line2);
nand2 M4_CalP1_SP4_SP9nc2_Xo3(M4_CalP1_SP4_SP9nc2_NotB, M4_CalP1_Propbus_4, M4_CalP1_SP4_SP9nc2_line3);
nand2 M4_CalP1_SP4_SP9nc2_Xo4(M4_CalP1_SP4_SP9nc2_line2, M4_CalP1_SP4_SP9nc2_line3, M4_CalP1_ParLo1);
inv M4_CalP1_SP5_SP7nc0_Xo0(M4_CalP1_Genbus_5, M4_CalP1_SP5_SP7nc0_NotA);
inv M4_CalP1_SP5_SP7nc0_Xo1(M4_CalP1_LocalC0_6, M4_CalP1_SP5_SP7nc0_NotB);
nand2 M4_CalP1_SP5_SP7nc0_Xo2(M4_CalP1_SP5_SP7nc0_NotA, M4_CalP1_LocalC0_6, M4_CalP1_SP5_SP7nc0_line2);
nand2 M4_CalP1_SP5_SP7nc0_Xo3(M4_CalP1_SP5_SP7nc0_NotB, M4_CalP1_Genbus_5, M4_CalP1_SP5_SP7nc0_line3);
nand2 M4_CalP1_SP5_SP7nc0_Xo4(M4_CalP1_SP5_SP7nc0_line2, M4_CalP1_SP5_SP7nc0_line3, M4_CalP1_SP5_line0);
inv M4_CalP1_SP5_SP7nc1_Xo0(M4_CalP1_LocalC0_7, M4_CalP1_SP5_SP7nc1_NotA);
inv M4_CalP1_SP5_SP7nc1_Xo1(M4_CalP1_SP5_line0, M4_CalP1_SP5_SP7nc1_NotB);
nand2 M4_CalP1_SP5_SP7nc1_Xo2(M4_CalP1_SP5_SP7nc1_NotA, M4_CalP1_SP5_line0, M4_CalP1_SP5_SP7nc1_line2);
nand2 M4_CalP1_SP5_SP7nc1_Xo3(M4_CalP1_SP5_SP7nc1_NotB, M4_CalP1_LocalC0_7, M4_CalP1_SP5_SP7nc1_line3);
nand2 M4_CalP1_SP5_SP7nc1_Xo4(M4_CalP1_SP5_SP7nc1_line2, M4_CalP1_SP5_SP7nc1_line3, M4_CalP1_SP5_line1);
inv M4_CalP1_SP5_SP7nc2_Xo0(M4_CalP1_Propbus_5, M4_CalP1_SP5_SP7nc2_NotA);
inv M4_CalP1_SP5_SP7nc2_Xo1(M4_CalP1_SP5_line1, M4_CalP1_SP5_SP7nc2_NotB);
nand2 M4_CalP1_SP5_SP7nc2_Xo2(M4_CalP1_SP5_SP7nc2_NotA, M4_CalP1_SP5_line1, M4_CalP1_SP5_SP7nc2_line2);
nand2 M4_CalP1_SP5_SP7nc2_Xo3(M4_CalP1_SP5_SP7nc2_NotB, M4_CalP1_Propbus_5, M4_CalP1_SP5_SP7nc2_line3);
nand2 M4_CalP1_SP5_SP7nc2_Xo4(M4_CalP1_SP5_SP7nc2_line2, M4_CalP1_SP5_SP7nc2_line3, M4_CalP1_SP5_line2);
inv M4_CalP1_SP5_SP7nc3_Xo0(M4_CalP1_Propbus_6, M4_CalP1_SP5_SP7nc3_NotA);
inv M4_CalP1_SP5_SP7nc3_Xo1(M4_CalP1_SP5_line2, M4_CalP1_SP5_SP7nc3_NotB);
nand2 M4_CalP1_SP5_SP7nc3_Xo2(M4_CalP1_SP5_SP7nc3_NotA, M4_CalP1_SP5_line2, M4_CalP1_SP5_SP7nc3_line2);
nand2 M4_CalP1_SP5_SP7nc3_Xo3(M4_CalP1_SP5_SP7nc3_NotB, M4_CalP1_Propbus_6, M4_CalP1_SP5_SP7nc3_line3);
nand2 M4_CalP1_SP5_SP7nc3_Xo4(M4_CalP1_SP5_SP7nc3_line2, M4_CalP1_SP5_SP7nc3_line3, M4_CalP1_SP5_line3);
inv M4_CalP1_SP5_SP7nc4_Xo0(M4_CalP1_Propbus_7, M4_CalP1_SP5_SP7nc4_NotA);
inv M4_CalP1_SP5_SP7nc4_Xo1(M4_CalP1_SP5_line3, M4_CalP1_SP5_SP7nc4_NotB);
nand2 M4_CalP1_SP5_SP7nc4_Xo2(M4_CalP1_SP5_SP7nc4_NotA, M4_CalP1_SP5_line3, M4_CalP1_SP5_SP7nc4_line2);
nand2 M4_CalP1_SP5_SP7nc4_Xo3(M4_CalP1_SP5_SP7nc4_NotB, M4_CalP1_Propbus_7, M4_CalP1_SP5_SP7nc4_line3);
nand2 M4_CalP1_SP5_SP7nc4_Xo4(M4_CalP1_SP5_SP7nc4_line2, M4_CalP1_SP5_SP7nc4_line3, M4_CalP1_SP5_line4);
inv M4_CalP1_SP5_SP7nc5_Xo0(M4_CalP1_Propbus_8, M4_CalP1_SP5_SP7nc5_NotA);
inv M4_CalP1_SP5_SP7nc5_Xo1(M4_CalP1_SP5_line4, M4_CalP1_SP5_SP7nc5_NotB);
nand2 M4_CalP1_SP5_SP7nc5_Xo2(M4_CalP1_SP5_SP7nc5_NotA, M4_CalP1_SP5_line4, M4_CalP1_SP5_SP7nc5_line2);
nand2 M4_CalP1_SP5_SP7nc5_Xo3(M4_CalP1_SP5_SP7nc5_NotB, M4_CalP1_Propbus_8, M4_CalP1_SP5_SP7nc5_line3);
nand2 M4_CalP1_SP5_SP7nc5_Xo4(M4_CalP1_SP5_SP7nc5_line2, M4_CalP1_SP5_SP7nc5_line3, M4_CalP1_ParHi0);
inv M4_CalP1_SP6_SP7c0(M4_CalP1_Propbus_8, M4_CalP1_SP6_NewInbus_6);
inv M4_CalP1_SP6_SP7c2_SP7nc0_Xo0(M4_CalP1_LocalC1_5, M4_CalP1_SP6_SP7c2_SP7nc0_NotA);
inv M4_CalP1_SP6_SP7c2_SP7nc0_Xo1(M4_CalP1_LocalC1_6, M4_CalP1_SP6_SP7c2_SP7nc0_NotB);
nand2 M4_CalP1_SP6_SP7c2_SP7nc0_Xo2(M4_CalP1_SP6_SP7c2_SP7nc0_NotA, M4_CalP1_LocalC1_6, M4_CalP1_SP6_SP7c2_SP7nc0_line2);
nand2 M4_CalP1_SP6_SP7c2_SP7nc0_Xo3(M4_CalP1_SP6_SP7c2_SP7nc0_NotB, M4_CalP1_LocalC1_5, M4_CalP1_SP6_SP7c2_SP7nc0_line3);
nand2 M4_CalP1_SP6_SP7c2_SP7nc0_Xo4(M4_CalP1_SP6_SP7c2_SP7nc0_line2, M4_CalP1_SP6_SP7c2_SP7nc0_line3, M4_CalP1_SP6_SP7c2_line0);
inv M4_CalP1_SP6_SP7c2_SP7nc1_Xo0(M4_CalP1_LocalC1_7, M4_CalP1_SP6_SP7c2_SP7nc1_NotA);
inv M4_CalP1_SP6_SP7c2_SP7nc1_Xo1(M4_CalP1_SP6_SP7c2_line0, M4_CalP1_SP6_SP7c2_SP7nc1_NotB);
nand2 M4_CalP1_SP6_SP7c2_SP7nc1_Xo2(M4_CalP1_SP6_SP7c2_SP7nc1_NotA, M4_CalP1_SP6_SP7c2_line0, M4_CalP1_SP6_SP7c2_SP7nc1_line2);
nand2 M4_CalP1_SP6_SP7c2_SP7nc1_Xo3(M4_CalP1_SP6_SP7c2_SP7nc1_NotB, M4_CalP1_LocalC1_7, M4_CalP1_SP6_SP7c2_SP7nc1_line3);
nand2 M4_CalP1_SP6_SP7c2_SP7nc1_Xo4(M4_CalP1_SP6_SP7c2_SP7nc1_line2, M4_CalP1_SP6_SP7c2_SP7nc1_line3, M4_CalP1_SP6_SP7c2_line1);
inv M4_CalP1_SP6_SP7c2_SP7nc2_Xo0(M4_CalP1_Propbus_5, M4_CalP1_SP6_SP7c2_SP7nc2_NotA);
inv M4_CalP1_SP6_SP7c2_SP7nc2_Xo1(M4_CalP1_SP6_SP7c2_line1, M4_CalP1_SP6_SP7c2_SP7nc2_NotB);
nand2 M4_CalP1_SP6_SP7c2_SP7nc2_Xo2(M4_CalP1_SP6_SP7c2_SP7nc2_NotA, M4_CalP1_SP6_SP7c2_line1, M4_CalP1_SP6_SP7c2_SP7nc2_line2);
nand2 M4_CalP1_SP6_SP7c2_SP7nc2_Xo3(M4_CalP1_SP6_SP7c2_SP7nc2_NotB, M4_CalP1_Propbus_5, M4_CalP1_SP6_SP7c2_SP7nc2_line3);
nand2 M4_CalP1_SP6_SP7c2_SP7nc2_Xo4(M4_CalP1_SP6_SP7c2_SP7nc2_line2, M4_CalP1_SP6_SP7c2_SP7nc2_line3, M4_CalP1_SP6_SP7c2_line2);
inv M4_CalP1_SP6_SP7c2_SP7nc3_Xo0(M4_CalP1_Propbus_6, M4_CalP1_SP6_SP7c2_SP7nc3_NotA);
inv M4_CalP1_SP6_SP7c2_SP7nc3_Xo1(M4_CalP1_SP6_SP7c2_line2, M4_CalP1_SP6_SP7c2_SP7nc3_NotB);
nand2 M4_CalP1_SP6_SP7c2_SP7nc3_Xo2(M4_CalP1_SP6_SP7c2_SP7nc3_NotA, M4_CalP1_SP6_SP7c2_line2, M4_CalP1_SP6_SP7c2_SP7nc3_line2);
nand2 M4_CalP1_SP6_SP7c2_SP7nc3_Xo3(M4_CalP1_SP6_SP7c2_SP7nc3_NotB, M4_CalP1_Propbus_6, M4_CalP1_SP6_SP7c2_SP7nc3_line3);
nand2 M4_CalP1_SP6_SP7c2_SP7nc3_Xo4(M4_CalP1_SP6_SP7c2_SP7nc3_line2, M4_CalP1_SP6_SP7c2_SP7nc3_line3, M4_CalP1_SP6_SP7c2_line3);
inv M4_CalP1_SP6_SP7c2_SP7nc4_Xo0(M4_CalP1_Propbus_7, M4_CalP1_SP6_SP7c2_SP7nc4_NotA);
inv M4_CalP1_SP6_SP7c2_SP7nc4_Xo1(M4_CalP1_SP6_SP7c2_line3, M4_CalP1_SP6_SP7c2_SP7nc4_NotB);
nand2 M4_CalP1_SP6_SP7c2_SP7nc4_Xo2(M4_CalP1_SP6_SP7c2_SP7nc4_NotA, M4_CalP1_SP6_SP7c2_line3, M4_CalP1_SP6_SP7c2_SP7nc4_line2);
nand2 M4_CalP1_SP6_SP7c2_SP7nc4_Xo3(M4_CalP1_SP6_SP7c2_SP7nc4_NotB, M4_CalP1_Propbus_7, M4_CalP1_SP6_SP7c2_SP7nc4_line3);
nand2 M4_CalP1_SP6_SP7c2_SP7nc4_Xo4(M4_CalP1_SP6_SP7c2_SP7nc4_line2, M4_CalP1_SP6_SP7c2_SP7nc4_line3, M4_CalP1_SP6_SP7c2_line4);
inv M4_CalP1_SP6_SP7c2_SP7nc5_Xo0(M4_CalP1_SP6_NewInbus_6, M4_CalP1_SP6_SP7c2_SP7nc5_NotA);
inv M4_CalP1_SP6_SP7c2_SP7nc5_Xo1(M4_CalP1_SP6_SP7c2_line4, M4_CalP1_SP6_SP7c2_SP7nc5_NotB);
nand2 M4_CalP1_SP6_SP7c2_SP7nc5_Xo2(M4_CalP1_SP6_SP7c2_SP7nc5_NotA, M4_CalP1_SP6_SP7c2_line4, M4_CalP1_SP6_SP7c2_SP7nc5_line2);
nand2 M4_CalP1_SP6_SP7c2_SP7nc5_Xo3(M4_CalP1_SP6_SP7c2_SP7nc5_NotB, M4_CalP1_SP6_NewInbus_6, M4_CalP1_SP6_SP7c2_SP7nc5_line3);
nand2 M4_CalP1_SP6_SP7c2_SP7nc5_Xo4(M4_CalP1_SP6_SP7c2_SP7nc5_line2, M4_CalP1_SP6_SP7c2_SP7nc5_line3, M4_CalP1_ParHi1);
inv M4_CalP1_SP7_Mux2_0(in1497, M4_CalP1_SP7_Not_ContIn);
and2 M4_CalP1_SP7_Mux2_1(M4_CalP1_ParLo0, M4_CalP1_SP7_Not_ContIn, M4_CalP1_SP7_line1);
and2 M4_CalP1_SP7_Mux2_2(M4_CalP1_ParLo1, in1497, M4_CalP1_SP7_line2);
or2 M4_CalP1_SP7_Mux2_3(M4_CalP1_SP7_line1, M4_CalP1_SP7_line2, M4_CalP1_ParLo);
inv M4_CalP1_SP8_Mux2_0(M4_CalP1_LocalC0_4, M4_CalP1_SP8_Not_ContIn);
and2 M4_CalP1_SP8_Mux2_1(M4_CalP1_ParHi0, M4_CalP1_SP8_Not_ContIn, M4_CalP1_SP8_line1);
and2 M4_CalP1_SP8_Mux2_2(M4_CalP1_ParHi1, M4_CalP1_LocalC0_4, M4_CalP1_SP8_line2);
or2 M4_CalP1_SP8_Mux2_3(M4_CalP1_SP8_line1, M4_CalP1_SP8_line2, M4_CalP1_ParHiCin0);
inv M4_CalP1_SP9_Mux2_0(M4_CalP1_LocalC1_4, M4_CalP1_SP9_Not_ContIn);
and2 M4_CalP1_SP9_Mux2_1(M4_CalP1_ParHi0, M4_CalP1_SP9_Not_ContIn, M4_CalP1_SP9_line1);
and2 M4_CalP1_SP9_Mux2_2(M4_CalP1_ParHi1, M4_CalP1_LocalC1_4, M4_CalP1_SP9_line2);
or2 M4_CalP1_SP9_Mux2_3(M4_CalP1_SP9_line1, M4_CalP1_SP9_line2, M4_CalP1_ParHiCin1);
inv M4_CalP1_SP10_Mux2_0(in1497, M4_CalP1_SP10_Not_ContIn);
and2 M4_CalP1_SP10_Mux2_1(M4_CalP1_ParHiCin0, M4_CalP1_SP10_Not_ContIn, M4_CalP1_SP10_line1);
and2 M4_CalP1_SP10_Mux2_2(M4_CalP1_ParHiCin1, in1497, M4_CalP1_SP10_line2);
or2 M4_CalP1_SP10_Mux2_3(M4_CalP1_SP10_line1, M4_CalP1_SP10_line2, M4_CalP1_ParHi);
inv M4_CalP1_SP11_Xo0(M4_CalP1_ParLo, M4_CalP1_SP11_NotA);
inv M4_CalP1_SP11_Xo1(M4_CalP1_ParHi, M4_CalP1_SP11_NotB);
nand2 M4_CalP1_SP11_Xo2(M4_CalP1_SP11_NotA, M4_CalP1_ParHi, M4_CalP1_SP11_line2);
nand2 M4_CalP1_SP11_Xo3(M4_CalP1_SP11_NotB, M4_CalP1_ParLo, M4_CalP1_SP11_line3);
nand2 M4_CalP1_SP11_Xo4(M4_CalP1_SP11_line2, M4_CalP1_SP11_line3, M4_SumPar);
inv M4_CalP2_M2M4_0(M4_LogicPar, M4_CalP2_NotLogicPar);
inv M4_CalP2_M2M4_1(M4_SumPar, M4_CalP2_NotSumPar);
inv M4_CalP2_M2M4_2_Mux2_0(in4091, M4_CalP2_M2M4_2_Not_ContIn);
and2 M4_CalP2_M2M4_2_Mux2_1(M4_CalP2_NotLogicPar, M4_CalP2_M2M4_2_Not_ContIn, M4_CalP2_M2M4_2_line1);
and2 M4_CalP2_M2M4_2_Mux2_2(M4_CalP2_NotSumPar, in4091, M4_CalP2_M2M4_2_line2);
or2 M4_CalP2_M2M4_2_Mux2_3(M4_CalP2_M2M4_2_line1, M4_CalP2_M2M4_2_line2, M4_CalP2_line0);
inv M4_CalP2_M2M4_3_Mux2_0(in4092, M4_CalP2_M2M4_3_Not_ContIn);
and2 M4_CalP2_M2M4_3_Mux2_1(M4_CalP2_line0, M4_CalP2_M2M4_3_Not_ContIn, M4_CalP2_M2M4_3_line1);
and2 M4_CalP2_M2M4_3_Mux2_2(in97, in4092, M4_CalP2_M2M4_3_line2);
or2 M4_CalP2_M2M4_3_Mux2_3(M4_CalP2_M2M4_3_line1, M4_CalP2_M2M4_3_line2, Not_SumLogicParY);
inv M4_CalP2_M2M4_4_Mux4_0(in4092, M4_CalP2_M2M4_4_Not_ContLo);
inv M4_CalP2_M2M4_4_Mux4_1(in4091, M4_CalP2_M2M4_4_Not_ContHi);
and3 M4_CalP2_M2M4_4_Mux4_2(M4_LogicPar, M4_CalP2_M2M4_4_Not_ContHi, M4_CalP2_M2M4_4_Not_ContLo, M4_CalP2_M2M4_4_line2);
and3 M4_CalP2_M2M4_4_Mux4_3(in118, M4_CalP2_M2M4_4_Not_ContHi, in4092, M4_CalP2_M2M4_4_line3);
and3 M4_CalP2_M2M4_4_Mux4_4(M4_SumPar, in4091, M4_CalP2_M2M4_4_Not_ContLo, M4_CalP2_M2M4_4_line4);
and3 M4_CalP2_M2M4_4_Mux4_5(vdd, in4091, in4092, M4_CalP2_M2M4_4_line5);
or4 M4_CalP2_M2M4_4_Mux4_6(M4_CalP2_M2M4_4_line2, M4_CalP2_M2M4_4_line3, M4_CalP2_M2M4_4_line4, M4_CalP2_M2M4_4_line5, out882);
inv M5_MP0_MXS0_Mux4_0(in1689, M5_MP0_MXS0_Not_ContLo);
inv M5_MP0_MXS0_Mux4_1(in1690, M5_MP0_MXS0_Not_ContHi);
and3 M5_MP0_MXS0_Mux4_2(Not_SumLogicParX, M5_MP0_MXS0_Not_ContHi, M5_MP0_MXS0_Not_ContLo, M5_MP0_MXS0_line2);
and3 M5_MP0_MXS0_Mux4_3(Not_SumLogicParY, M5_MP0_MXS0_Not_ContHi, in1689, M5_MP0_MXS0_line3);
and3 M5_MP0_MXS0_Mux4_4(in176, in1690, M5_MP0_MXS0_Not_ContLo, M5_MP0_MXS0_line4);
and3 M5_MP0_MXS0_Mux4_5(in179, in1690, in1689, M5_MP0_MXS0_line5);
or4 M5_MP0_MXS0_Mux4_6(M5_MP0_MXS0_line2, M5_MP0_MXS0_line3, M5_MP0_MXS0_line4, M5_MP0_MXS0_line5, M5_MP0_tempOut1);
inv M5_MP0_MXS1_Mux4_0(in1691, M5_MP0_MXS1_Not_ContLo);
inv M5_MP0_MXS1_Mux4_1(in1694, M5_MP0_MXS1_Not_ContHi);
and3 M5_MP0_MXS1_Mux4_2(Not_SumLogicParX, M5_MP0_MXS1_Not_ContHi, M5_MP0_MXS1_Not_ContLo, M5_MP0_MXS1_line2);
and3 M5_MP0_MXS1_Mux4_3(Not_SumLogicParY, M5_MP0_MXS1_Not_ContHi, in1691, M5_MP0_MXS1_line3);
and3 M5_MP0_MXS1_Mux4_4(in176, in1694, M5_MP0_MXS1_Not_ContLo, M5_MP0_MXS1_line4);
and3 M5_MP0_MXS1_Mux4_5(in179, in1694, in1691, M5_MP0_MXS1_line5);
or4 M5_MP0_MXS1_Mux4_6(M5_MP0_MXS1_line2, M5_MP0_MXS1_line3, M5_MP0_MXS1_line4, M5_MP0_MXS1_line5, M5_MP0_tempOut2);
inv M5_MP0_MXS2_Mux4_0(in4088, M5_MP0_MXS2_Not_ContLo);
inv M5_MP0_MXS2_Mux4_1(in4087, M5_MP0_MXS2_Not_ContHi);
and3 M5_MP0_MXS2_Mux4_2(Not_SumLogicParX, M5_MP0_MXS2_Not_ContHi, M5_MP0_MXS2_Not_ContLo, M5_MP0_MXS2_line2);
and3 M5_MP0_MXS2_Mux4_3(Not_SumLogicParY, M5_MP0_MXS2_Not_ContHi, in4088, M5_MP0_MXS2_line3);
and3 M5_MP0_MXS2_Mux4_4(in14, in4087, M5_MP0_MXS2_Not_ContLo, M5_MP0_MXS2_line4);
and3 M5_MP0_MXS2_Mux4_5(in64, in4087, in4088, M5_MP0_MXS2_line5);
or4 M5_MP0_MXS2_Mux4_6(M5_MP0_MXS2_line2, M5_MP0_MXS2_line3, M5_MP0_MXS2_line4, M5_MP0_MXS2_line5, out767);
inv M5_MP0_MXS3_Mux4_0(in4089, M5_MP0_MXS3_Not_ContLo);
inv M5_MP0_MXS3_Mux4_1(in4090, M5_MP0_MXS3_Not_ContHi);
and3 M5_MP0_MXS3_Mux4_2(Not_SumLogicParX, M5_MP0_MXS3_Not_ContHi, M5_MP0_MXS3_Not_ContLo, M5_MP0_MXS3_line2);
and3 M5_MP0_MXS3_Mux4_3(Not_SumLogicParY, M5_MP0_MXS3_Not_ContHi, in4089, M5_MP0_MXS3_line3);
and3 M5_MP0_MXS3_Mux4_4(in14, in4090, M5_MP0_MXS3_Not_ContLo, M5_MP0_MXS3_line4);
and3 M5_MP0_MXS3_Mux4_5(in64, in4090, in4089, M5_MP0_MXS3_line5);
or4 M5_MP0_MXS3_Mux4_6(M5_MP0_MXS3_line2, M5_MP0_MXS3_line3, M5_MP0_MXS3_line4, M5_MP0_MXS3_line5, out807);
and2 M5_MP0_MXS4(M5_MP0_tempOut1, in137, M5_NotOP1);
and2 M5_MP0_MXS5(M5_MP0_tempOut2, in137, M5_NotOP2);
inv M5_MP1(M5_NotOP1, out658);
inv M5_MP2(M5_NotOP2, out690);
inv M0_Inv4_0(in3548, NotContLogic3_0_0);
inv M0_Inv4_1(in3546, NotContLogic3_0_1);
inv M0_Inv4_2(in3550, NotContLogic3_0_2);
inv M0_Inv4_3(in3552, NotContLogic3_0_3);
inv M6_CSL0_CL0_LB0_Mux2_0(in361, M6_CSL0_CL0_LB0_Not_ContIn);
and2 M6_CSL0_CL0_LB0_Mux2_1(in254, M6_CSL0_CL0_LB0_Not_ContIn, M6_CSL0_CL0_LB0_line1);
and2 M6_CSL0_CL0_LB0_Mux2_2(in242, in361, M6_CSL0_CL0_LB0_line2);
or2 M6_CSL0_CL0_LB0_Mux2_3(M6_CSL0_CL0_LB0_line1, M6_CSL0_CL0_LB0_line2, M6_CSL0_CL0_line0);
inv M6_CSL0_CL0_LB1_Mux2_0(in361, M6_CSL0_CL0_LB1_Not_ContIn);
and2 M6_CSL0_CL0_LB1_Mux2_1(in251, M6_CSL0_CL0_LB1_Not_ContIn, M6_CSL0_CL0_LB1_line1);
and2 M6_CSL0_CL0_LB1_Mux2_2(in248, in361, M6_CSL0_CL0_LB1_line2);
or2 M6_CSL0_CL0_LB1_Mux2_3(M6_CSL0_CL0_LB1_line1, M6_CSL0_CL0_LB1_line2, M6_CSL0_CL0_line1);
or2 M6_CSL0_CL0_LB2(vdd, M6_CSL0_CL0_line0, M6_CSL0_CL0_line2);
nand2 M6_CSL0_CL0_LB3(vdd, M6_CSL0_CL0_line1, M6_CSL0_CL0_line3);
and2 M6_CSL0_CL0_LB4(M6_CSL0_CL0_line2, M6_CSL0_CL0_line3, LogicXbus_0);
inv M6_CSL0_CL1_LB0_Mux2_0(in351, M6_CSL0_CL1_LB0_Not_ContIn);
and2 M6_CSL0_CL1_LB0_Mux2_1(NotContLogic3_0_0, M6_CSL0_CL1_LB0_Not_ContIn, M6_CSL0_CL1_LB0_line1);
and2 M6_CSL0_CL1_LB0_Mux2_2(NotContLogic3_0_1, in351, M6_CSL0_CL1_LB0_line2);
or2 M6_CSL0_CL1_LB0_Mux2_3(M6_CSL0_CL1_LB0_line1, M6_CSL0_CL1_LB0_line2, M6_CSL0_CL1_line0);
inv M6_CSL0_CL1_LB1_Mux2_0(in351, M6_CSL0_CL1_LB1_Not_ContIn);
and2 M6_CSL0_CL1_LB1_Mux2_1(NotContLogic3_0_2, M6_CSL0_CL1_LB1_Not_ContIn, M6_CSL0_CL1_LB1_line1);
and2 M6_CSL0_CL1_LB1_Mux2_2(NotContLogic3_0_3, in351, M6_CSL0_CL1_LB1_line2);
or2 M6_CSL0_CL1_LB1_Mux2_3(M6_CSL0_CL1_LB1_line1, M6_CSL0_CL1_LB1_line2, M6_CSL0_CL1_line1);
or2 M6_CSL0_CL1_LB2(in534, M6_CSL0_CL1_line0, M6_CSL0_CL1_line2);
nand2 M6_CSL0_CL1_LB3(in534, M6_CSL0_CL1_line1, M6_CSL0_CL1_line3);
and2 M6_CSL0_CL1_LB4(M6_CSL0_CL1_line2, M6_CSL0_CL1_line3, LogicXbus_1);
inv M6_CSL0_CL2_LB0_Mux2_0(in341, M6_CSL0_CL2_LB0_Not_ContIn);
and2 M6_CSL0_CL2_LB0_Mux2_1(NotContLogic3_0_0, M6_CSL0_CL2_LB0_Not_ContIn, M6_CSL0_CL2_LB0_line1);
and2 M6_CSL0_CL2_LB0_Mux2_2(NotContLogic3_0_1, in341, M6_CSL0_CL2_LB0_line2);
or2 M6_CSL0_CL2_LB0_Mux2_3(M6_CSL0_CL2_LB0_line1, M6_CSL0_CL2_LB0_line2, M6_CSL0_CL2_line0);
inv M6_CSL0_CL2_LB1_Mux2_0(in341, M6_CSL0_CL2_LB1_Not_ContIn);
and2 M6_CSL0_CL2_LB1_Mux2_1(NotContLogic3_0_2, M6_CSL0_CL2_LB1_Not_ContIn, M6_CSL0_CL2_LB1_line1);
and2 M6_CSL0_CL2_LB1_Mux2_2(NotContLogic3_0_3, in341, M6_CSL0_CL2_LB1_line2);
or2 M6_CSL0_CL2_LB1_Mux2_3(M6_CSL0_CL2_LB1_line1, M6_CSL0_CL2_LB1_line2, M6_CSL0_CL2_line1);
or2 M6_CSL0_CL2_LB2(in523, M6_CSL0_CL2_line0, M6_CSL0_CL2_line2);
nand2 M6_CSL0_CL2_LB3(in523, M6_CSL0_CL2_line1, M6_CSL0_CL2_line3);
and2 M6_CSL0_CL2_LB4(M6_CSL0_CL2_line2, M6_CSL0_CL2_line3, LogicXbus_2);
inv M6_CSL0_CL3_LB0_Mux2_0(vdd, M6_CSL0_CL3_LB0_Not_ContIn);
and2 M6_CSL0_CL3_LB0_Mux2_1(NotContLogic3_0_0, M6_CSL0_CL3_LB0_Not_ContIn, M6_CSL0_CL3_LB0_line1);
and2 M6_CSL0_CL3_LB0_Mux2_2(NotContLogic3_0_1, vdd, M6_CSL0_CL3_LB0_line2);
or2 M6_CSL0_CL3_LB0_Mux2_3(M6_CSL0_CL3_LB0_line1, M6_CSL0_CL3_LB0_line2, M6_CSL0_CL3_line0);
inv M6_CSL0_CL3_LB1_Mux2_0(vdd, M6_CSL0_CL3_LB1_Not_ContIn);
and2 M6_CSL0_CL3_LB1_Mux2_1(NotContLogic3_0_2, M6_CSL0_CL3_LB1_Not_ContIn, M6_CSL0_CL3_LB1_line1);
and2 M6_CSL0_CL3_LB1_Mux2_2(NotContLogic3_0_3, vdd, M6_CSL0_CL3_LB1_line2);
or2 M6_CSL0_CL3_LB1_Mux2_3(M6_CSL0_CL3_LB1_line1, M6_CSL0_CL3_LB1_line2, M6_CSL0_CL3_line1);
or2 M6_CSL0_CL3_LB2(in514, M6_CSL0_CL3_line0, M6_CSL0_CL3_line2);
nand2 M6_CSL0_CL3_LB3(in514, M6_CSL0_CL3_line1, M6_CSL0_CL3_line3);
and2 M6_CSL0_CL3_LB4(M6_CSL0_CL3_line2, M6_CSL0_CL3_line3, LogicXbus_3);
inv M6_CSL0_CL4_LB0_Mux2_0(in324, M6_CSL0_CL4_LB0_Not_ContIn);
and2 M6_CSL0_CL4_LB0_Mux2_1(NotContLogic3_0_0, M6_CSL0_CL4_LB0_Not_ContIn, M6_CSL0_CL4_LB0_line1);
and2 M6_CSL0_CL4_LB0_Mux2_2(NotContLogic3_0_1, in324, M6_CSL0_CL4_LB0_line2);
or2 M6_CSL0_CL4_LB0_Mux2_3(M6_CSL0_CL4_LB0_line1, M6_CSL0_CL4_LB0_line2, M6_CSL0_CL4_line0);
inv M6_CSL0_CL4_LB1_Mux2_0(in324, M6_CSL0_CL4_LB1_Not_ContIn);
and2 M6_CSL0_CL4_LB1_Mux2_1(NotContLogic3_0_2, M6_CSL0_CL4_LB1_Not_ContIn, M6_CSL0_CL4_LB1_line1);
and2 M6_CSL0_CL4_LB1_Mux2_2(NotContLogic3_0_3, in324, M6_CSL0_CL4_LB1_line2);
or2 M6_CSL0_CL4_LB1_Mux2_3(M6_CSL0_CL4_LB1_line1, M6_CSL0_CL4_LB1_line2, M6_CSL0_CL4_line1);
or2 M6_CSL0_CL4_LB2(in503, M6_CSL0_CL4_line0, M6_CSL0_CL4_line2);
nand2 M6_CSL0_CL4_LB3(in503, M6_CSL0_CL4_line1, M6_CSL0_CL4_line3);
and2 M6_CSL0_CL4_LB4(M6_CSL0_CL4_line2, M6_CSL0_CL4_line3, LogicXbus_4);
inv M6_CSL0_CL5_LB0_Mux2_0(in316, M6_CSL0_CL5_LB0_Not_ContIn);
and2 M6_CSL0_CL5_LB0_Mux2_1(in254, M6_CSL0_CL5_LB0_Not_ContIn, M6_CSL0_CL5_LB0_line1);
and2 M6_CSL0_CL5_LB0_Mux2_2(in242, in316, M6_CSL0_CL5_LB0_line2);
or2 M6_CSL0_CL5_LB0_Mux2_3(M6_CSL0_CL5_LB0_line1, M6_CSL0_CL5_LB0_line2, M6_CSL0_CL5_line0);
inv M6_CSL0_CL5_LB1_Mux2_0(in316, M6_CSL0_CL5_LB1_Not_ContIn);
and2 M6_CSL0_CL5_LB1_Mux2_1(in251, M6_CSL0_CL5_LB1_Not_ContIn, M6_CSL0_CL5_LB1_line1);
and2 M6_CSL0_CL5_LB1_Mux2_2(in248, in316, M6_CSL0_CL5_LB1_line2);
or2 M6_CSL0_CL5_LB1_Mux2_3(M6_CSL0_CL5_LB1_line1, M6_CSL0_CL5_LB1_line2, M6_CSL0_CL5_line1);
or2 M6_CSL0_CL5_LB2(in490, M6_CSL0_CL5_line0, M6_CSL0_CL5_line2);
nand2 M6_CSL0_CL5_LB3(in490, M6_CSL0_CL5_line1, M6_CSL0_CL5_line3);
and2 M6_CSL0_CL5_LB4(M6_CSL0_CL5_line2, M6_CSL0_CL5_line3, LogicXbus_5);
inv M6_CSL0_CL6_LB0_Mux2_0(in308, M6_CSL0_CL6_LB0_Not_ContIn);
and2 M6_CSL0_CL6_LB0_Mux2_1(in254, M6_CSL0_CL6_LB0_Not_ContIn, M6_CSL0_CL6_LB0_line1);
and2 M6_CSL0_CL6_LB0_Mux2_2(in242, in308, M6_CSL0_CL6_LB0_line2);
or2 M6_CSL0_CL6_LB0_Mux2_3(M6_CSL0_CL6_LB0_line1, M6_CSL0_CL6_LB0_line2, M6_CSL0_CL6_line0);
inv M6_CSL0_CL6_LB1_Mux2_0(in308, M6_CSL0_CL6_LB1_Not_ContIn);
and2 M6_CSL0_CL6_LB1_Mux2_1(in251, M6_CSL0_CL6_LB1_Not_ContIn, M6_CSL0_CL6_LB1_line1);
and2 M6_CSL0_CL6_LB1_Mux2_2(in248, in308, M6_CSL0_CL6_LB1_line2);
or2 M6_CSL0_CL6_LB1_Mux2_3(M6_CSL0_CL6_LB1_line1, M6_CSL0_CL6_LB1_line2, M6_CSL0_CL6_line1);
or2 M6_CSL0_CL6_LB2(in479, M6_CSL0_CL6_line0, M6_CSL0_CL6_line2);
nand2 M6_CSL0_CL6_LB3(in479, M6_CSL0_CL6_line1, M6_CSL0_CL6_line3);
and2 M6_CSL0_CL6_LB4(M6_CSL0_CL6_line2, M6_CSL0_CL6_line3, LogicXbus_6);
inv M6_CSL0_CL7_LB0_Mux2_0(in302, M6_CSL0_CL7_LB0_Not_ContIn);
and2 M6_CSL0_CL7_LB0_Mux2_1(in254, M6_CSL0_CL7_LB0_Not_ContIn, M6_CSL0_CL7_LB0_line1);
and2 M6_CSL0_CL7_LB0_Mux2_2(in242, in302, M6_CSL0_CL7_LB0_line2);
or2 M6_CSL0_CL7_LB0_Mux2_3(M6_CSL0_CL7_LB0_line1, M6_CSL0_CL7_LB0_line2, M6_CSL0_CL7_line0);
inv M6_CSL0_CL7_LB1_Mux2_0(in302, M6_CSL0_CL7_LB1_Not_ContIn);
and2 M6_CSL0_CL7_LB1_Mux2_1(in251, M6_CSL0_CL7_LB1_Not_ContIn, M6_CSL0_CL7_LB1_line1);
and2 M6_CSL0_CL7_LB1_Mux2_2(in248, in302, M6_CSL0_CL7_LB1_line2);
or2 M6_CSL0_CL7_LB1_Mux2_3(M6_CSL0_CL7_LB1_line1, M6_CSL0_CL7_LB1_line2, M6_CSL0_CL7_line1);
or2 M6_CSL0_CL7_LB2(vdd, M6_CSL0_CL7_line0, M6_CSL0_CL7_line2);
nand2 M6_CSL0_CL7_LB3(vdd, M6_CSL0_CL7_line1, M6_CSL0_CL7_line3);
and2 M6_CSL0_CL7_LB4(M6_CSL0_CL7_line2, M6_CSL0_CL7_line3, LogicXbus_7);
inv M6_CSL0_CL8_LB0_Mux2_0(in293, M6_CSL0_CL8_LB0_Not_ContIn);
and2 M6_CSL0_CL8_LB0_Mux2_1(in254, M6_CSL0_CL8_LB0_Not_ContIn, M6_CSL0_CL8_LB0_line1);
and2 M6_CSL0_CL8_LB0_Mux2_2(in242, in293, M6_CSL0_CL8_LB0_line2);
or2 M6_CSL0_CL8_LB0_Mux2_3(M6_CSL0_CL8_LB0_line1, M6_CSL0_CL8_LB0_line2, M6_CSL0_CL8_line0);
inv M6_CSL0_CL8_LB1_Mux2_0(in293, M6_CSL0_CL8_LB1_Not_ContIn);
and2 M6_CSL0_CL8_LB1_Mux2_1(in251, M6_CSL0_CL8_LB1_Not_ContIn, M6_CSL0_CL8_LB1_line1);
and2 M6_CSL0_CL8_LB1_Mux2_2(in248, in293, M6_CSL0_CL8_LB1_line2);
or2 M6_CSL0_CL8_LB1_Mux2_3(M6_CSL0_CL8_LB1_line1, M6_CSL0_CL8_LB1_line2, M6_CSL0_CL8_line1);
or2 M6_CSL0_CL8_LB2(gnd, M6_CSL0_CL8_line0, M6_CSL0_CL8_line2);
nand2 M6_CSL0_CL8_LB3(gnd, M6_CSL0_CL8_line1, M6_CSL0_CL8_line3);
and2 M6_CSL0_CL8_LB4(M6_CSL0_CL8_line2, M6_CSL0_CL8_line3, LogicXbus_8);
and2 M6_CSL1_Add0_GP9_0(Xbus_0, vdd, M6_CSL1_Genbus_0);
and2 M6_CSL1_Add0_GP9_1(Xbus_1, in534, M6_CSL1_Genbus_1);
and2 M6_CSL1_Add0_GP9_2(Xbus_2, in523, M6_CSL1_Genbus_2);
and2 M6_CSL1_Add0_GP9_3(Xbus_3, in514, M6_CSL1_Genbus_3);
and2 M6_CSL1_Add0_GP9_4(Xbus_4, in503, M6_CSL1_Genbus_4);
and2 M6_CSL1_Add0_GP9_5(Xbus_5, in490, M6_CSL1_Genbus_5);
and2 M6_CSL1_Add0_GP9_6(Xbus_6, in479, M6_CSL1_Genbus_6);
and2 M6_CSL1_Add0_GP9_7(Xbus_7, vdd, M6_CSL1_Genbus_7);
and2 M6_CSL1_Add0_GP9_8(Xbus_8, vdd, M6_CSL1_Genbus_8);
inv M6_CSL1_Add0_GP9_9_Xo0(Xbus_0, M6_CSL1_Add0_GP9_9_NotA);
inv M6_CSL1_Add0_GP9_9_Xo1(vdd, M6_CSL1_Add0_GP9_9_NotB);
nand2 M6_CSL1_Add0_GP9_9_Xo2(M6_CSL1_Add0_GP9_9_NotA, vdd, M6_CSL1_Add0_GP9_9_line2);
nand2 M6_CSL1_Add0_GP9_9_Xo3(M6_CSL1_Add0_GP9_9_NotB, Xbus_0, M6_CSL1_Add0_GP9_9_line3);
nand2 M6_CSL1_Add0_GP9_9_Xo4(M6_CSL1_Add0_GP9_9_line2, M6_CSL1_Add0_GP9_9_line3, M6_CSL1_Propbus_0);
inv M6_CSL1_Add0_GP9_10_Xo0(Xbus_1, M6_CSL1_Add0_GP9_10_NotA);
inv M6_CSL1_Add0_GP9_10_Xo1(in534, M6_CSL1_Add0_GP9_10_NotB);
nand2 M6_CSL1_Add0_GP9_10_Xo2(M6_CSL1_Add0_GP9_10_NotA, in534, M6_CSL1_Add0_GP9_10_line2);
nand2 M6_CSL1_Add0_GP9_10_Xo3(M6_CSL1_Add0_GP9_10_NotB, Xbus_1, M6_CSL1_Add0_GP9_10_line3);
nand2 M6_CSL1_Add0_GP9_10_Xo4(M6_CSL1_Add0_GP9_10_line2, M6_CSL1_Add0_GP9_10_line3, M6_CSL1_Propbus_1);
inv M6_CSL1_Add0_GP9_11_Xo0(Xbus_2, M6_CSL1_Add0_GP9_11_NotA);
inv M6_CSL1_Add0_GP9_11_Xo1(in523, M6_CSL1_Add0_GP9_11_NotB);
nand2 M6_CSL1_Add0_GP9_11_Xo2(M6_CSL1_Add0_GP9_11_NotA, in523, M6_CSL1_Add0_GP9_11_line2);
nand2 M6_CSL1_Add0_GP9_11_Xo3(M6_CSL1_Add0_GP9_11_NotB, Xbus_2, M6_CSL1_Add0_GP9_11_line3);
nand2 M6_CSL1_Add0_GP9_11_Xo4(M6_CSL1_Add0_GP9_11_line2, M6_CSL1_Add0_GP9_11_line3, M6_CSL1_Propbus_2);
inv M6_CSL1_Add0_GP9_12_Xo0(Xbus_3, M6_CSL1_Add0_GP9_12_NotA);
inv M6_CSL1_Add0_GP9_12_Xo1(in514, M6_CSL1_Add0_GP9_12_NotB);
nand2 M6_CSL1_Add0_GP9_12_Xo2(M6_CSL1_Add0_GP9_12_NotA, in514, M6_CSL1_Add0_GP9_12_line2);
nand2 M6_CSL1_Add0_GP9_12_Xo3(M6_CSL1_Add0_GP9_12_NotB, Xbus_3, M6_CSL1_Add0_GP9_12_line3);
nand2 M6_CSL1_Add0_GP9_12_Xo4(M6_CSL1_Add0_GP9_12_line2, M6_CSL1_Add0_GP9_12_line3, M6_CSL1_Propbus_3);
inv M6_CSL1_Add0_GP9_13_Xo0(Xbus_4, M6_CSL1_Add0_GP9_13_NotA);
inv M6_CSL1_Add0_GP9_13_Xo1(in503, M6_CSL1_Add0_GP9_13_NotB);
nand2 M6_CSL1_Add0_GP9_13_Xo2(M6_CSL1_Add0_GP9_13_NotA, in503, M6_CSL1_Add0_GP9_13_line2);
nand2 M6_CSL1_Add0_GP9_13_Xo3(M6_CSL1_Add0_GP9_13_NotB, Xbus_4, M6_CSL1_Add0_GP9_13_line3);
nand2 M6_CSL1_Add0_GP9_13_Xo4(M6_CSL1_Add0_GP9_13_line2, M6_CSL1_Add0_GP9_13_line3, M6_CSL1_Propbus_4);
inv M6_CSL1_Add0_GP9_14_Xo0(Xbus_5, M6_CSL1_Add0_GP9_14_NotA);
inv M6_CSL1_Add0_GP9_14_Xo1(in490, M6_CSL1_Add0_GP9_14_NotB);
nand2 M6_CSL1_Add0_GP9_14_Xo2(M6_CSL1_Add0_GP9_14_NotA, in490, M6_CSL1_Add0_GP9_14_line2);
nand2 M6_CSL1_Add0_GP9_14_Xo3(M6_CSL1_Add0_GP9_14_NotB, Xbus_5, M6_CSL1_Add0_GP9_14_line3);
nand2 M6_CSL1_Add0_GP9_14_Xo4(M6_CSL1_Add0_GP9_14_line2, M6_CSL1_Add0_GP9_14_line3, M6_CSL1_Propbus_5);
inv M6_CSL1_Add0_GP9_15_Xo0(Xbus_6, M6_CSL1_Add0_GP9_15_NotA);
inv M6_CSL1_Add0_GP9_15_Xo1(in479, M6_CSL1_Add0_GP9_15_NotB);
nand2 M6_CSL1_Add0_GP9_15_Xo2(M6_CSL1_Add0_GP9_15_NotA, in479, M6_CSL1_Add0_GP9_15_line2);
nand2 M6_CSL1_Add0_GP9_15_Xo3(M6_CSL1_Add0_GP9_15_NotB, Xbus_6, M6_CSL1_Add0_GP9_15_line3);
nand2 M6_CSL1_Add0_GP9_15_Xo4(M6_CSL1_Add0_GP9_15_line2, M6_CSL1_Add0_GP9_15_line3, M6_CSL1_Propbus_6);
inv M6_CSL1_Add0_GP9_16_Xo0(Xbus_7, M6_CSL1_Add0_GP9_16_NotA);
inv M6_CSL1_Add0_GP9_16_Xo1(vdd, M6_CSL1_Add0_GP9_16_NotB);
nand2 M6_CSL1_Add0_GP9_16_Xo2(M6_CSL1_Add0_GP9_16_NotA, vdd, M6_CSL1_Add0_GP9_16_line2);
nand2 M6_CSL1_Add0_GP9_16_Xo3(M6_CSL1_Add0_GP9_16_NotB, Xbus_7, M6_CSL1_Add0_GP9_16_line3);
nand2 M6_CSL1_Add0_GP9_16_Xo4(M6_CSL1_Add0_GP9_16_line2, M6_CSL1_Add0_GP9_16_line3, M6_CSL1_Propbus_7);
inv M6_CSL1_Add0_GP9_17_Xo0(Xbus_8, M6_CSL1_Add0_GP9_17_NotA);
inv M6_CSL1_Add0_GP9_17_Xo1(vdd, M6_CSL1_Add0_GP9_17_NotB);
nand2 M6_CSL1_Add0_GP9_17_Xo2(M6_CSL1_Add0_GP9_17_NotA, vdd, M6_CSL1_Add0_GP9_17_line2);
nand2 M6_CSL1_Add0_GP9_17_Xo3(M6_CSL1_Add0_GP9_17_NotB, Xbus_8, M6_CSL1_Add0_GP9_17_line3);
nand2 M6_CSL1_Add0_GP9_17_Xo4(M6_CSL1_Add0_GP9_17_line2, M6_CSL1_Add0_GP9_17_line3, M6_CSL1_Propbus_8);
and2 M6_CSL1_Add1_CB0_Ao2_0(M6_CSL1_Propbus_0, in54, M6_CSL1_Add1_CB0_line0);
or2 M6_CSL1_Add1_CB0_Ao2_1(M6_CSL1_Genbus_0, M6_CSL1_Add1_CB0_line0, M6_CSL1_Carry_0);
and2 M6_CSL1_Add1_CB1_Ao3a_0(M6_CSL1_Propbus_1, M6_CSL1_Genbus_0, M6_CSL1_Add1_CB1_line0);
and3 M6_CSL1_Add1_CB1_Ao3a_1(M6_CSL1_Propbus_1, M6_CSL1_Propbus_0, in54, M6_CSL1_Add1_CB1_line1);
or3 M6_CSL1_Add1_CB1_Ao3a_2(M6_CSL1_Genbus_1, M6_CSL1_Add1_CB1_line0, M6_CSL1_Add1_CB1_line1, M6_CSL1_Carry_1);
and2 M6_CSL1_Add1_CB2_Ao4a_0(M6_CSL1_Propbus_2, M6_CSL1_Genbus_1, M6_CSL1_Add1_CB2_line0);
and3 M6_CSL1_Add1_CB2_Ao4a_1(M6_CSL1_Propbus_2, M6_CSL1_Propbus_1, M6_CSL1_Genbus_0, M6_CSL1_Add1_CB2_line1);
and4 M6_CSL1_Add1_CB2_Ao4a_2(M6_CSL1_Propbus_2, M6_CSL1_Propbus_1, M6_CSL1_Propbus_0, in54, M6_CSL1_Add1_CB2_line2);
or4 M6_CSL1_Add1_CB2_Ao4a_3(M6_CSL1_Genbus_2, M6_CSL1_Add1_CB2_line0, M6_CSL1_Add1_CB2_line1, M6_CSL1_Add1_CB2_line2, M6_CSL1_Carry_2);
and2 M6_CSL1_Add1_CB3_Ao5a_0(M6_CSL1_Propbus_3, M6_CSL1_Genbus_2, M6_CSL1_Add1_CB3_line0);
and3 M6_CSL1_Add1_CB3_Ao5a_1(M6_CSL1_Propbus_3, M6_CSL1_Propbus_2, M6_CSL1_Genbus_1, M6_CSL1_Add1_CB3_line1);
and4 M6_CSL1_Add1_CB3_Ao5a_2(M6_CSL1_Propbus_3, M6_CSL1_Propbus_2, M6_CSL1_Propbus_1, M6_CSL1_Genbus_0, M6_CSL1_Add1_CB3_line2);
and5 M6_CSL1_Add1_CB3_Ao5a_3(M6_CSL1_Propbus_3, M6_CSL1_Propbus_2, M6_CSL1_Propbus_1, M6_CSL1_Propbus_0, in54, M6_CSL1_Add1_CB3_line3);
or5 M6_CSL1_Add1_CB3_Ao5a_4(M6_CSL1_Genbus_3, M6_CSL1_Add1_CB3_line0, M6_CSL1_Add1_CB3_line1, M6_CSL1_Add1_CB3_line2, M6_CSL1_Add1_CB3_line3, M6_CSL1_Carry_3);
and2 M6_CSL1_Add1_CB4_Ao5a_0(M6_CSL1_Propbus_4, M6_CSL1_Genbus_3, M6_CSL1_Add1_CB4_line0);
and3 M6_CSL1_Add1_CB4_Ao5a_1(M6_CSL1_Propbus_4, M6_CSL1_Propbus_3, M6_CSL1_Genbus_2, M6_CSL1_Add1_CB4_line1);
and4 M6_CSL1_Add1_CB4_Ao5a_2(M6_CSL1_Propbus_4, M6_CSL1_Propbus_3, M6_CSL1_Propbus_2, M6_CSL1_Genbus_1, M6_CSL1_Add1_CB4_line2);
and5 M6_CSL1_Add1_CB4_Ao5a_3(M6_CSL1_Propbus_4, M6_CSL1_Propbus_3, M6_CSL1_Propbus_2, M6_CSL1_Propbus_1, M6_CSL1_Genbus_0, M6_CSL1_Add1_CB4_line3);
or5 M6_CSL1_Add1_CB4_Ao5a_4(M6_CSL1_Genbus_4, M6_CSL1_Add1_CB4_line0, M6_CSL1_Add1_CB4_line1, M6_CSL1_Add1_CB4_line2, M6_CSL1_Add1_CB4_line3, M6_CSL1_Add1_LocalC0_4);
and5 M6_CSL1_Add1_CB5(M6_CSL1_Propbus_0, M6_CSL1_Propbus_1, M6_CSL1_Propbus_2, M6_CSL1_Propbus_3, M6_CSL1_Propbus_4, M6_CSL1_Add1_Prop4_0);
and2 M6_CSL1_Add1_CB6(in54, M6_CSL1_Add1_Prop4_0, M6_CSL1_Add1_PropCin);
or2 M6_CSL1_Add1_CB7(M6_CSL1_Add1_LocalC0_4, M6_CSL1_Add1_PropCin, M6_CSL1_Carry_4);
and2 M6_CSL1_Add1_CB8_Ao5a_0(M6_CSL1_Propbus_8, M6_CSL1_Genbus_7, M6_CSL1_Add1_CB8_line0);
and3 M6_CSL1_Add1_CB8_Ao5a_1(M6_CSL1_Propbus_8, M6_CSL1_Propbus_7, M6_CSL1_Genbus_6, M6_CSL1_Add1_CB8_line1);
and4 M6_CSL1_Add1_CB8_Ao5a_2(M6_CSL1_Propbus_8, M6_CSL1_Propbus_7, M6_CSL1_Propbus_6, M6_CSL1_Genbus_5, M6_CSL1_Add1_CB8_line2);
and5 M6_CSL1_Add1_CB8_Ao5a_3(M6_CSL1_Propbus_8, M6_CSL1_Propbus_7, M6_CSL1_Propbus_6, M6_CSL1_Propbus_5, M6_CSL1_Add1_LocalC0_4, M6_CSL1_Add1_CB8_line3);
or5 M6_CSL1_Add1_CB8_Ao5a_4(M6_CSL1_Genbus_8, M6_CSL1_Add1_CB8_line0, M6_CSL1_Add1_CB8_line1, M6_CSL1_Add1_CB8_line2, M6_CSL1_Add1_CB8_line3, out629);
and4 M6_CSL1_Add1_CB9(M6_CSL1_Propbus_5, M6_CSL1_Propbus_6, M6_CSL1_Propbus_7, M6_CSL1_Propbus_8, M6_CSL1_Add1_Prop8_5);
and2 M6_CSL1_Add1_CB10(M6_CSL1_Add1_Prop4_0, M6_CSL1_Add1_Prop8_5, out615);
or2 M6_CSL1_Add2_GLC4_0(M6_CSL1_Genbus_5, M6_CSL1_Propbus_5, M6_CSL1_LocalHC1_0);
and2 M6_CSL1_Add2_GLC4_1_Ao2_0(M6_CSL1_Propbus_6, M6_CSL1_Genbus_5, M6_CSL1_Add2_GLC4_1_line0);
or2 M6_CSL1_Add2_GLC4_1_Ao2_1(M6_CSL1_Genbus_6, M6_CSL1_Add2_GLC4_1_line0, M6_CSL1_LocalHC0_1);
and2 M6_CSL1_Add2_GLC4_2_Ao3a_0(M6_CSL1_Propbus_6, M6_CSL1_Genbus_5, M6_CSL1_Add2_GLC4_2_line0);
and2 M6_CSL1_Add2_GLC4_2_Ao3a_1(M6_CSL1_Propbus_6, M6_CSL1_Propbus_5, M6_CSL1_Add2_GLC4_2_line1);
or3 M6_CSL1_Add2_GLC4_2_Ao3a_2(M6_CSL1_Genbus_6, M6_CSL1_Add2_GLC4_2_line0, M6_CSL1_Add2_GLC4_2_line1, M6_CSL1_LocalHC1_1);
and2 M6_CSL1_Add2_GLC4_3_Ao3a_0(M6_CSL1_Propbus_7, M6_CSL1_Genbus_6, M6_CSL1_Add2_GLC4_3_line0);
and3 M6_CSL1_Add2_GLC4_3_Ao3a_1(M6_CSL1_Propbus_7, M6_CSL1_Propbus_6, M6_CSL1_Genbus_5, M6_CSL1_Add2_GLC4_3_line1);
or3 M6_CSL1_Add2_GLC4_3_Ao3a_2(M6_CSL1_Genbus_7, M6_CSL1_Add2_GLC4_3_line0, M6_CSL1_Add2_GLC4_3_line1, M6_CSL1_LocalHC0_2);
and2 M6_CSL1_Add2_GLC4_4_Ao4a_0(M6_CSL1_Propbus_7, M6_CSL1_Genbus_6, M6_CSL1_Add2_GLC4_4_line0);
and3 M6_CSL1_Add2_GLC4_4_Ao4a_1(M6_CSL1_Propbus_7, M6_CSL1_Propbus_6, M6_CSL1_Genbus_5, M6_CSL1_Add2_GLC4_4_line1);
and3 M6_CSL1_Add2_GLC4_4_Ao4a_2(M6_CSL1_Propbus_7, M6_CSL1_Propbus_6, M6_CSL1_Propbus_5, M6_CSL1_Add2_GLC4_4_line2);
or4 M6_CSL1_Add2_GLC4_4_Ao4a_3(M6_CSL1_Genbus_7, M6_CSL1_Add2_GLC4_4_line0, M6_CSL1_Add2_GLC4_4_line1, M6_CSL1_Add2_GLC4_4_line2, M6_CSL1_LocalHC1_2);
inv M6_CSL1_Add3_X2a6_0_Xo0(M6_CSL1_Propbus_0, M6_CSL1_Add3_X2a6_0_NotA);
inv M6_CSL1_Add3_X2a6_0_Xo1(in54, M6_CSL1_Add3_X2a6_0_NotB);
nand2 M6_CSL1_Add3_X2a6_0_Xo2(M6_CSL1_Add3_X2a6_0_NotA, in54, M6_CSL1_Add3_X2a6_0_line2);
nand2 M6_CSL1_Add3_X2a6_0_Xo3(M6_CSL1_Add3_X2a6_0_NotB, M6_CSL1_Propbus_0, M6_CSL1_Add3_X2a6_0_line3);
nand2 M6_CSL1_Add3_X2a6_0_Xo4(M6_CSL1_Add3_X2a6_0_line2, M6_CSL1_Add3_X2a6_0_line3, SumXbus_0);
inv M6_CSL1_Add3_X2a6_1_Xo0(M6_CSL1_Propbus_1, M6_CSL1_Add3_X2a6_1_NotA);
inv M6_CSL1_Add3_X2a6_1_Xo1(M6_CSL1_Carry_0, M6_CSL1_Add3_X2a6_1_NotB);
nand2 M6_CSL1_Add3_X2a6_1_Xo2(M6_CSL1_Add3_X2a6_1_NotA, M6_CSL1_Carry_0, M6_CSL1_Add3_X2a6_1_line2);
nand2 M6_CSL1_Add3_X2a6_1_Xo3(M6_CSL1_Add3_X2a6_1_NotB, M6_CSL1_Propbus_1, M6_CSL1_Add3_X2a6_1_line3);
nand2 M6_CSL1_Add3_X2a6_1_Xo4(M6_CSL1_Add3_X2a6_1_line2, M6_CSL1_Add3_X2a6_1_line3, SumXbus_1);
inv M6_CSL1_Add3_X2a6_2_Xo0(M6_CSL1_Propbus_2, M6_CSL1_Add3_X2a6_2_NotA);
inv M6_CSL1_Add3_X2a6_2_Xo1(M6_CSL1_Carry_1, M6_CSL1_Add3_X2a6_2_NotB);
nand2 M6_CSL1_Add3_X2a6_2_Xo2(M6_CSL1_Add3_X2a6_2_NotA, M6_CSL1_Carry_1, M6_CSL1_Add3_X2a6_2_line2);
nand2 M6_CSL1_Add3_X2a6_2_Xo3(M6_CSL1_Add3_X2a6_2_NotB, M6_CSL1_Propbus_2, M6_CSL1_Add3_X2a6_2_line3);
nand2 M6_CSL1_Add3_X2a6_2_Xo4(M6_CSL1_Add3_X2a6_2_line2, M6_CSL1_Add3_X2a6_2_line3, SumXbus_2);
inv M6_CSL1_Add3_X2a6_3_Xo0(M6_CSL1_Propbus_3, M6_CSL1_Add3_X2a6_3_NotA);
inv M6_CSL1_Add3_X2a6_3_Xo1(M6_CSL1_Carry_2, M6_CSL1_Add3_X2a6_3_NotB);
nand2 M6_CSL1_Add3_X2a6_3_Xo2(M6_CSL1_Add3_X2a6_3_NotA, M6_CSL1_Carry_2, M6_CSL1_Add3_X2a6_3_line2);
nand2 M6_CSL1_Add3_X2a6_3_Xo3(M6_CSL1_Add3_X2a6_3_NotB, M6_CSL1_Propbus_3, M6_CSL1_Add3_X2a6_3_line3);
nand2 M6_CSL1_Add3_X2a6_3_Xo4(M6_CSL1_Add3_X2a6_3_line2, M6_CSL1_Add3_X2a6_3_line3, SumXbus_3);
inv M6_CSL1_Add3_X2a6_4_Xo0(M6_CSL1_Propbus_4, M6_CSL1_Add3_X2a6_4_NotA);
inv M6_CSL1_Add3_X2a6_4_Xo1(M6_CSL1_Carry_3, M6_CSL1_Add3_X2a6_4_NotB);
nand2 M6_CSL1_Add3_X2a6_4_Xo2(M6_CSL1_Add3_X2a6_4_NotA, M6_CSL1_Carry_3, M6_CSL1_Add3_X2a6_4_line2);
nand2 M6_CSL1_Add3_X2a6_4_Xo3(M6_CSL1_Add3_X2a6_4_NotB, M6_CSL1_Propbus_4, M6_CSL1_Add3_X2a6_4_line3);
nand2 M6_CSL1_Add3_X2a6_4_Xo4(M6_CSL1_Add3_X2a6_4_line2, M6_CSL1_Add3_X2a6_4_line3, SumXbus_4);
inv M6_CSL1_Add3_X2a6_5_Xo0(M6_CSL1_Propbus_5, M6_CSL1_Add3_X2a6_5_NotA);
inv M6_CSL1_Add3_X2a6_5_Xo1(M6_CSL1_Carry_4, M6_CSL1_Add3_X2a6_5_NotB);
nand2 M6_CSL1_Add3_X2a6_5_Xo2(M6_CSL1_Add3_X2a6_5_NotA, M6_CSL1_Carry_4, M6_CSL1_Add3_X2a6_5_line2);
nand2 M6_CSL1_Add3_X2a6_5_Xo3(M6_CSL1_Add3_X2a6_5_NotB, M6_CSL1_Propbus_5, M6_CSL1_Add3_X2a6_5_line3);
nand2 M6_CSL1_Add3_X2a6_5_Xo4(M6_CSL1_Add3_X2a6_5_line2, M6_CSL1_Add3_X2a6_5_line3, SumXbus_5);
inv M6_CSL1_Add4_X2a6_0_Xo0(M6_CSL1_Propbus_6, M6_CSL1_Add4_X2a6_0_NotA);
inv M6_CSL1_Add4_X2a6_0_Xo1(M6_CSL1_Genbus_5, M6_CSL1_Add4_X2a6_0_NotB);
nand2 M6_CSL1_Add4_X2a6_0_Xo2(M6_CSL1_Add4_X2a6_0_NotA, M6_CSL1_Genbus_5, M6_CSL1_Add4_X2a6_0_line2);
nand2 M6_CSL1_Add4_X2a6_0_Xo3(M6_CSL1_Add4_X2a6_0_NotB, M6_CSL1_Propbus_6, M6_CSL1_Add4_X2a6_0_line3);
nand2 M6_CSL1_Add4_X2a6_0_Xo4(M6_CSL1_Add4_X2a6_0_line2, M6_CSL1_Add4_X2a6_0_line3, M6_CSL1_SumH01bus_0);
inv M6_CSL1_Add4_X2a6_1_Xo0(M6_CSL1_Propbus_7, M6_CSL1_Add4_X2a6_1_NotA);
inv M6_CSL1_Add4_X2a6_1_Xo1(M6_CSL1_LocalHC0_1, M6_CSL1_Add4_X2a6_1_NotB);
nand2 M6_CSL1_Add4_X2a6_1_Xo2(M6_CSL1_Add4_X2a6_1_NotA, M6_CSL1_LocalHC0_1, M6_CSL1_Add4_X2a6_1_line2);
nand2 M6_CSL1_Add4_X2a6_1_Xo3(M6_CSL1_Add4_X2a6_1_NotB, M6_CSL1_Propbus_7, M6_CSL1_Add4_X2a6_1_line3);
nand2 M6_CSL1_Add4_X2a6_1_Xo4(M6_CSL1_Add4_X2a6_1_line2, M6_CSL1_Add4_X2a6_1_line3, M6_CSL1_SumH01bus_1);
inv M6_CSL1_Add4_X2a6_2_Xo0(M6_CSL1_Propbus_8, M6_CSL1_Add4_X2a6_2_NotA);
inv M6_CSL1_Add4_X2a6_2_Xo1(M6_CSL1_LocalHC0_2, M6_CSL1_Add4_X2a6_2_NotB);
nand2 M6_CSL1_Add4_X2a6_2_Xo2(M6_CSL1_Add4_X2a6_2_NotA, M6_CSL1_LocalHC0_2, M6_CSL1_Add4_X2a6_2_line2);
nand2 M6_CSL1_Add4_X2a6_2_Xo3(M6_CSL1_Add4_X2a6_2_NotB, M6_CSL1_Propbus_8, M6_CSL1_Add4_X2a6_2_line3);
nand2 M6_CSL1_Add4_X2a6_2_Xo4(M6_CSL1_Add4_X2a6_2_line2, M6_CSL1_Add4_X2a6_2_line3, M6_CSL1_SumH01bus_2);
inv M6_CSL1_Add4_X2a6_3_Xo0(M6_CSL1_Propbus_6, M6_CSL1_Add4_X2a6_3_NotA);
inv M6_CSL1_Add4_X2a6_3_Xo1(M6_CSL1_LocalHC1_0, M6_CSL1_Add4_X2a6_3_NotB);
nand2 M6_CSL1_Add4_X2a6_3_Xo2(M6_CSL1_Add4_X2a6_3_NotA, M6_CSL1_LocalHC1_0, M6_CSL1_Add4_X2a6_3_line2);
nand2 M6_CSL1_Add4_X2a6_3_Xo3(M6_CSL1_Add4_X2a6_3_NotB, M6_CSL1_Propbus_6, M6_CSL1_Add4_X2a6_3_line3);
nand2 M6_CSL1_Add4_X2a6_3_Xo4(M6_CSL1_Add4_X2a6_3_line2, M6_CSL1_Add4_X2a6_3_line3, M6_CSL1_SumH01bus_3);
inv M6_CSL1_Add4_X2a6_4_Xo0(M6_CSL1_Propbus_7, M6_CSL1_Add4_X2a6_4_NotA);
inv M6_CSL1_Add4_X2a6_4_Xo1(M6_CSL1_LocalHC1_1, M6_CSL1_Add4_X2a6_4_NotB);
nand2 M6_CSL1_Add4_X2a6_4_Xo2(M6_CSL1_Add4_X2a6_4_NotA, M6_CSL1_LocalHC1_1, M6_CSL1_Add4_X2a6_4_line2);
nand2 M6_CSL1_Add4_X2a6_4_Xo3(M6_CSL1_Add4_X2a6_4_NotB, M6_CSL1_Propbus_7, M6_CSL1_Add4_X2a6_4_line3);
nand2 M6_CSL1_Add4_X2a6_4_Xo4(M6_CSL1_Add4_X2a6_4_line2, M6_CSL1_Add4_X2a6_4_line3, M6_CSL1_SumH01bus_4);
inv M6_CSL1_Add4_X2a6_5_Xo0(M6_CSL1_Propbus_8, M6_CSL1_Add4_X2a6_5_NotA);
inv M6_CSL1_Add4_X2a6_5_Xo1(M6_CSL1_LocalHC1_2, M6_CSL1_Add4_X2a6_5_NotB);
nand2 M6_CSL1_Add4_X2a6_5_Xo2(M6_CSL1_Add4_X2a6_5_NotA, M6_CSL1_LocalHC1_2, M6_CSL1_Add4_X2a6_5_line2);
nand2 M6_CSL1_Add4_X2a6_5_Xo3(M6_CSL1_Add4_X2a6_5_NotB, M6_CSL1_Propbus_8, M6_CSL1_Add4_X2a6_5_line3);
nand2 M6_CSL1_Add4_X2a6_5_Xo4(M6_CSL1_Add4_X2a6_5_line2, M6_CSL1_Add4_X2a6_5_line3, M6_CSL1_SumH01bus_5);
inv M6_CSL1_Add5_Mux2_0(M6_CSL1_Carry_4, M6_CSL1_Add5_Not_ContIn);
and2 M6_CSL1_Add5_Mux2_1(M6_CSL1_SumH01bus_0, M6_CSL1_Add5_Not_ContIn, M6_CSL1_Add5_line1);
and2 M6_CSL1_Add5_Mux2_2(M6_CSL1_SumH01bus_3, M6_CSL1_Carry_4, M6_CSL1_Add5_line2);
or2 M6_CSL1_Add5_Mux2_3(M6_CSL1_Add5_line1, M6_CSL1_Add5_line2, SumXbus_6);
inv M6_CSL1_Add6_Mux2_0(M6_CSL1_Carry_4, M6_CSL1_Add6_Not_ContIn);
and2 M6_CSL1_Add6_Mux2_1(M6_CSL1_SumH01bus_1, M6_CSL1_Add6_Not_ContIn, M6_CSL1_Add6_line1);
and2 M6_CSL1_Add6_Mux2_2(M6_CSL1_SumH01bus_4, M6_CSL1_Carry_4, M6_CSL1_Add6_line2);
or2 M6_CSL1_Add6_Mux2_3(M6_CSL1_Add6_line1, M6_CSL1_Add6_line2, SumXbus_7);
inv M6_CSL1_Add7_Mux2_0(M6_CSL1_Carry_4, M6_CSL1_Add7_Not_ContIn);
and2 M6_CSL1_Add7_Mux2_1(M6_CSL1_SumH01bus_2, M6_CSL1_Add7_Not_ContIn, M6_CSL1_Add7_line1);
and2 M6_CSL1_Add7_Mux2_2(M6_CSL1_SumH01bus_5, M6_CSL1_Carry_4, M6_CSL1_Add7_line2);
or2 M6_CSL1_Add7_Mux2_3(M6_CSL1_Add7_line1, M6_CSL1_Add7_line2, SumXbus_8);
inv M6_CSL2_Mx9_0_Mx4_0_Mux4_0(in4092, M6_CSL2_Mx9_0_Mx4_0_Not_ContLo);
inv M6_CSL2_Mx9_0_Mx4_0_Mux4_1(in4091, M6_CSL2_Mx9_0_Mx4_0_Not_ContHi);
and3 M6_CSL2_Mx9_0_Mx4_0_Mux4_2(LogicXbus_0, M6_CSL2_Mx9_0_Mx4_0_Not_ContHi, M6_CSL2_Mx9_0_Mx4_0_Not_ContLo, M6_CSL2_Mx9_0_Mx4_0_line2);
and3 M6_CSL2_Mx9_0_Mx4_0_Mux4_3(in131, M6_CSL2_Mx9_0_Mx4_0_Not_ContHi, in4092, M6_CSL2_Mx9_0_Mx4_0_line3);
and3 M6_CSL2_Mx9_0_Mx4_0_Mux4_4(SumXbus_0, in4091, M6_CSL2_Mx9_0_Mx4_0_Not_ContLo, M6_CSL2_Mx9_0_Mx4_0_line4);
and3 M6_CSL2_Mx9_0_Mx4_0_Mux4_5(gnd, in4091, in4092, M6_CSL2_Mx9_0_Mx4_0_line5);
or4 M6_CSL2_Mx9_0_Mx4_0_Mux4_6(M6_CSL2_Mx9_0_Mx4_0_line2, M6_CSL2_Mx9_0_Mx4_0_line3, M6_CSL2_Mx9_0_Mx4_0_line4, M6_CSL2_Mx9_0_Mx4_0_line5, FXbus_0);
inv M6_CSL2_Mx9_0_Mx4_1_Mux4_0(in4092, M6_CSL2_Mx9_0_Mx4_1_Not_ContLo);
inv M6_CSL2_Mx9_0_Mx4_1_Mux4_1(in4091, M6_CSL2_Mx9_0_Mx4_1_Not_ContHi);
and3 M6_CSL2_Mx9_0_Mx4_1_Mux4_2(LogicXbus_1, M6_CSL2_Mx9_0_Mx4_1_Not_ContHi, M6_CSL2_Mx9_0_Mx4_1_Not_ContLo, M6_CSL2_Mx9_0_Mx4_1_line2);
and3 M6_CSL2_Mx9_0_Mx4_1_Mux4_3(in129, M6_CSL2_Mx9_0_Mx4_1_Not_ContHi, in4092, M6_CSL2_Mx9_0_Mx4_1_line3);
and3 M6_CSL2_Mx9_0_Mx4_1_Mux4_4(SumXbus_1, in4091, M6_CSL2_Mx9_0_Mx4_1_Not_ContLo, M6_CSL2_Mx9_0_Mx4_1_line4);
and3 M6_CSL2_Mx9_0_Mx4_1_Mux4_5(gnd, in4091, in4092, M6_CSL2_Mx9_0_Mx4_1_line5);
or4 M6_CSL2_Mx9_0_Mx4_1_Mux4_6(M6_CSL2_Mx9_0_Mx4_1_line2, M6_CSL2_Mx9_0_Mx4_1_line3, M6_CSL2_Mx9_0_Mx4_1_line4, M6_CSL2_Mx9_0_Mx4_1_line5, FXbus_1);
inv M6_CSL2_Mx9_0_Mx4_2_Mux4_0(in4092, M6_CSL2_Mx9_0_Mx4_2_Not_ContLo);
inv M6_CSL2_Mx9_0_Mx4_2_Mux4_1(in4091, M6_CSL2_Mx9_0_Mx4_2_Not_ContHi);
and3 M6_CSL2_Mx9_0_Mx4_2_Mux4_2(LogicXbus_2, M6_CSL2_Mx9_0_Mx4_2_Not_ContHi, M6_CSL2_Mx9_0_Mx4_2_Not_ContLo, M6_CSL2_Mx9_0_Mx4_2_line2);
and3 M6_CSL2_Mx9_0_Mx4_2_Mux4_3(in119, M6_CSL2_Mx9_0_Mx4_2_Not_ContHi, in4092, M6_CSL2_Mx9_0_Mx4_2_line3);
and3 M6_CSL2_Mx9_0_Mx4_2_Mux4_4(SumXbus_2, in4091, M6_CSL2_Mx9_0_Mx4_2_Not_ContLo, M6_CSL2_Mx9_0_Mx4_2_line4);
and3 M6_CSL2_Mx9_0_Mx4_2_Mux4_5(gnd, in4091, in4092, M6_CSL2_Mx9_0_Mx4_2_line5);
or4 M6_CSL2_Mx9_0_Mx4_2_Mux4_6(M6_CSL2_Mx9_0_Mx4_2_line2, M6_CSL2_Mx9_0_Mx4_2_line3, M6_CSL2_Mx9_0_Mx4_2_line4, M6_CSL2_Mx9_0_Mx4_2_line5, FXbus_2);
inv M6_CSL2_Mx9_0_Mx4_3_Mux4_0(in4092, M6_CSL2_Mx9_0_Mx4_3_Not_ContLo);
inv M6_CSL2_Mx9_0_Mx4_3_Mux4_1(in4091, M6_CSL2_Mx9_0_Mx4_3_Not_ContHi);
and3 M6_CSL2_Mx9_0_Mx4_3_Mux4_2(LogicXbus_3, M6_CSL2_Mx9_0_Mx4_3_Not_ContHi, M6_CSL2_Mx9_0_Mx4_3_Not_ContLo, M6_CSL2_Mx9_0_Mx4_3_line2);
and3 M6_CSL2_Mx9_0_Mx4_3_Mux4_3(in130, M6_CSL2_Mx9_0_Mx4_3_Not_ContHi, in4092, M6_CSL2_Mx9_0_Mx4_3_line3);
and3 M6_CSL2_Mx9_0_Mx4_3_Mux4_4(SumXbus_3, in4091, M6_CSL2_Mx9_0_Mx4_3_Not_ContLo, M6_CSL2_Mx9_0_Mx4_3_line4);
and3 M6_CSL2_Mx9_0_Mx4_3_Mux4_5(gnd, in4091, in4092, M6_CSL2_Mx9_0_Mx4_3_line5);
or4 M6_CSL2_Mx9_0_Mx4_3_Mux4_6(M6_CSL2_Mx9_0_Mx4_3_line2, M6_CSL2_Mx9_0_Mx4_3_line3, M6_CSL2_Mx9_0_Mx4_3_line4, M6_CSL2_Mx9_0_Mx4_3_line5, FXbus_3);
inv M6_CSL2_Mx9_1_Mx4_0_Mux4_0(in4092, M6_CSL2_Mx9_1_Mx4_0_Not_ContLo);
inv M6_CSL2_Mx9_1_Mx4_0_Mux4_1(in4091, M6_CSL2_Mx9_1_Mx4_0_Not_ContHi);
and3 M6_CSL2_Mx9_1_Mx4_0_Mux4_2(LogicXbus_4, M6_CSL2_Mx9_1_Mx4_0_Not_ContHi, M6_CSL2_Mx9_1_Mx4_0_Not_ContLo, M6_CSL2_Mx9_1_Mx4_0_line2);
and3 M6_CSL2_Mx9_1_Mx4_0_Mux4_3(in52, M6_CSL2_Mx9_1_Mx4_0_Not_ContHi, in4092, M6_CSL2_Mx9_1_Mx4_0_line3);
and3 M6_CSL2_Mx9_1_Mx4_0_Mux4_4(SumXbus_4, in4091, M6_CSL2_Mx9_1_Mx4_0_Not_ContLo, M6_CSL2_Mx9_1_Mx4_0_line4);
and3 M6_CSL2_Mx9_1_Mx4_0_Mux4_5(gnd, in4091, in4092, M6_CSL2_Mx9_1_Mx4_0_line5);
or4 M6_CSL2_Mx9_1_Mx4_0_Mux4_6(M6_CSL2_Mx9_1_Mx4_0_line2, M6_CSL2_Mx9_1_Mx4_0_line3, M6_CSL2_Mx9_1_Mx4_0_line4, M6_CSL2_Mx9_1_Mx4_0_line5, FXbus_4);
inv M6_CSL2_Mx9_1_Mx4_1_Mux4_0(in4092, M6_CSL2_Mx9_1_Mx4_1_Not_ContLo);
inv M6_CSL2_Mx9_1_Mx4_1_Mux4_1(in4091, M6_CSL2_Mx9_1_Mx4_1_Not_ContHi);
and3 M6_CSL2_Mx9_1_Mx4_1_Mux4_2(LogicXbus_5, M6_CSL2_Mx9_1_Mx4_1_Not_ContHi, M6_CSL2_Mx9_1_Mx4_1_Not_ContLo, M6_CSL2_Mx9_1_Mx4_1_line2);
and3 M6_CSL2_Mx9_1_Mx4_1_Mux4_3(in112, M6_CSL2_Mx9_1_Mx4_1_Not_ContHi, in4092, M6_CSL2_Mx9_1_Mx4_1_line3);
and3 M6_CSL2_Mx9_1_Mx4_1_Mux4_4(SumXbus_5, in4091, M6_CSL2_Mx9_1_Mx4_1_Not_ContLo, M6_CSL2_Mx9_1_Mx4_1_line4);
and3 M6_CSL2_Mx9_1_Mx4_1_Mux4_5(gnd, in4091, in4092, M6_CSL2_Mx9_1_Mx4_1_line5);
or4 M6_CSL2_Mx9_1_Mx4_1_Mux4_6(M6_CSL2_Mx9_1_Mx4_1_line2, M6_CSL2_Mx9_1_Mx4_1_line3, M6_CSL2_Mx9_1_Mx4_1_line4, M6_CSL2_Mx9_1_Mx4_1_line5, FXbus_5);
inv M6_CSL2_Mx9_1_Mx4_2_Mux4_0(in4092, M6_CSL2_Mx9_1_Mx4_2_Not_ContLo);
inv M6_CSL2_Mx9_1_Mx4_2_Mux4_1(in4091, M6_CSL2_Mx9_1_Mx4_2_Not_ContHi);
and3 M6_CSL2_Mx9_1_Mx4_2_Mux4_2(LogicXbus_6, M6_CSL2_Mx9_1_Mx4_2_Not_ContHi, M6_CSL2_Mx9_1_Mx4_2_Not_ContLo, M6_CSL2_Mx9_1_Mx4_2_line2);
and3 M6_CSL2_Mx9_1_Mx4_2_Mux4_3(in116, M6_CSL2_Mx9_1_Mx4_2_Not_ContHi, in4092, M6_CSL2_Mx9_1_Mx4_2_line3);
and3 M6_CSL2_Mx9_1_Mx4_2_Mux4_4(SumXbus_6, in4091, M6_CSL2_Mx9_1_Mx4_2_Not_ContLo, M6_CSL2_Mx9_1_Mx4_2_line4);
and3 M6_CSL2_Mx9_1_Mx4_2_Mux4_5(gnd, in4091, in4092, M6_CSL2_Mx9_1_Mx4_2_line5);
or4 M6_CSL2_Mx9_1_Mx4_2_Mux4_6(M6_CSL2_Mx9_1_Mx4_2_line2, M6_CSL2_Mx9_1_Mx4_2_line3, M6_CSL2_Mx9_1_Mx4_2_line4, M6_CSL2_Mx9_1_Mx4_2_line5, FXbus_6);
inv M6_CSL2_Mx9_1_Mx4_3_Mux4_0(in4092, M6_CSL2_Mx9_1_Mx4_3_Not_ContLo);
inv M6_CSL2_Mx9_1_Mx4_3_Mux4_1(in4091, M6_CSL2_Mx9_1_Mx4_3_Not_ContHi);
and3 M6_CSL2_Mx9_1_Mx4_3_Mux4_2(LogicXbus_7, M6_CSL2_Mx9_1_Mx4_3_Not_ContHi, M6_CSL2_Mx9_1_Mx4_3_Not_ContLo, M6_CSL2_Mx9_1_Mx4_3_line2);
and3 M6_CSL2_Mx9_1_Mx4_3_Mux4_3(in121, M6_CSL2_Mx9_1_Mx4_3_Not_ContHi, in4092, M6_CSL2_Mx9_1_Mx4_3_line3);
and3 M6_CSL2_Mx9_1_Mx4_3_Mux4_4(SumXbus_7, in4091, M6_CSL2_Mx9_1_Mx4_3_Not_ContLo, M6_CSL2_Mx9_1_Mx4_3_line4);
and3 M6_CSL2_Mx9_1_Mx4_3_Mux4_5(gnd, in4091, in4092, M6_CSL2_Mx9_1_Mx4_3_line5);
or4 M6_CSL2_Mx9_1_Mx4_3_Mux4_6(M6_CSL2_Mx9_1_Mx4_3_line2, M6_CSL2_Mx9_1_Mx4_3_line3, M6_CSL2_Mx9_1_Mx4_3_line4, M6_CSL2_Mx9_1_Mx4_3_line5, FXbus_7);
inv M6_CSL2_Mx9_2_Mux4_0(in4092, M6_CSL2_Mx9_2_Not_ContLo);
inv M6_CSL2_Mx9_2_Mux4_1(in4091, M6_CSL2_Mx9_2_Not_ContHi);
and3 M6_CSL2_Mx9_2_Mux4_2(LogicXbus_8, M6_CSL2_Mx9_2_Not_ContHi, M6_CSL2_Mx9_2_Not_ContLo, M6_CSL2_Mx9_2_line2);
and3 M6_CSL2_Mx9_2_Mux4_3(in123, M6_CSL2_Mx9_2_Not_ContHi, in4092, M6_CSL2_Mx9_2_line3);
and3 M6_CSL2_Mx9_2_Mux4_4(SumXbus_8, in4091, M6_CSL2_Mx9_2_Not_ContLo, M6_CSL2_Mx9_2_line4);
and3 M6_CSL2_Mx9_2_Mux4_5(gnd, in4091, in4092, M6_CSL2_Mx9_2_line5);
or4 M6_CSL2_Mx9_2_Mux4_6(M6_CSL2_Mx9_2_line2, M6_CSL2_Mx9_2_line3, M6_CSL2_Mx9_2_line4, M6_CSL2_Mx9_2_line5, FXbus_8);
inv M7_CSL0_CL0_LB0_Mux2_0(in281, M7_CSL0_CL0_LB0_Not_ContIn);
and2 M7_CSL0_CL0_LB0_Mux2_1(NotContLogic3_0_0, M7_CSL0_CL0_LB0_Not_ContIn, M7_CSL0_CL0_LB0_line1);
and2 M7_CSL0_CL0_LB0_Mux2_2(NotContLogic3_0_1, in281, M7_CSL0_CL0_LB0_line2);
or2 M7_CSL0_CL0_LB0_Mux2_3(M7_CSL0_CL0_LB0_line1, M7_CSL0_CL0_LB0_line2, M7_CSL0_CL0_line0);
inv M7_CSL0_CL0_LB1_Mux2_0(in281, M7_CSL0_CL0_LB1_Not_ContIn);
and2 M7_CSL0_CL0_LB1_Mux2_1(NotContLogic3_0_2, M7_CSL0_CL0_LB1_Not_ContIn, M7_CSL0_CL0_LB1_line1);
and2 M7_CSL0_CL0_LB1_Mux2_2(NotContLogic3_0_3, in281, M7_CSL0_CL0_LB1_line2);
or2 M7_CSL0_CL0_LB1_Mux2_3(M7_CSL0_CL0_LB1_line1, M7_CSL0_CL0_LB1_line2, M7_CSL0_CL0_line1);
or2 M7_CSL0_CL0_LB2(in374, M7_CSL0_CL0_line0, M7_CSL0_CL0_line2);
nand2 M7_CSL0_CL0_LB3(in374, M7_CSL0_CL0_line1, M7_CSL0_CL0_line3);
and2 M7_CSL0_CL0_LB4(M7_CSL0_CL0_line2, M7_CSL0_CL0_line3, LogicYbus_0);
inv M7_CSL0_CL1_LB0_Mux2_0(in273, M7_CSL0_CL1_LB0_Not_ContIn);
and2 M7_CSL0_CL1_LB0_Mux2_1(NotContLogic3_0_0, M7_CSL0_CL1_LB0_Not_ContIn, M7_CSL0_CL1_LB0_line1);
and2 M7_CSL0_CL1_LB0_Mux2_2(NotContLogic3_0_1, in273, M7_CSL0_CL1_LB0_line2);
or2 M7_CSL0_CL1_LB0_Mux2_3(M7_CSL0_CL1_LB0_line1, M7_CSL0_CL1_LB0_line2, M7_CSL0_CL1_line0);
inv M7_CSL0_CL1_LB1_Mux2_0(in273, M7_CSL0_CL1_LB1_Not_ContIn);
and2 M7_CSL0_CL1_LB1_Mux2_1(NotContLogic3_0_2, M7_CSL0_CL1_LB1_Not_ContIn, M7_CSL0_CL1_LB1_line1);
and2 M7_CSL0_CL1_LB1_Mux2_2(NotContLogic3_0_3, in273, M7_CSL0_CL1_LB1_line2);
or2 M7_CSL0_CL1_LB1_Mux2_3(M7_CSL0_CL1_LB1_line1, M7_CSL0_CL1_LB1_line2, M7_CSL0_CL1_line1);
or2 M7_CSL0_CL1_LB2(in411, M7_CSL0_CL1_line0, M7_CSL0_CL1_line2);
nand2 M7_CSL0_CL1_LB3(in411, M7_CSL0_CL1_line1, M7_CSL0_CL1_line3);
and2 M7_CSL0_CL1_LB4(M7_CSL0_CL1_line2, M7_CSL0_CL1_line3, LogicYbus_1);
inv M7_CSL0_CL2_LB0_Mux2_0(in265, M7_CSL0_CL2_LB0_Not_ContIn);
and2 M7_CSL0_CL2_LB0_Mux2_1(NotContLogic3_0_0, M7_CSL0_CL2_LB0_Not_ContIn, M7_CSL0_CL2_LB0_line1);
and2 M7_CSL0_CL2_LB0_Mux2_2(NotContLogic3_0_1, in265, M7_CSL0_CL2_LB0_line2);
or2 M7_CSL0_CL2_LB0_Mux2_3(M7_CSL0_CL2_LB0_line1, M7_CSL0_CL2_LB0_line2, M7_CSL0_CL2_line0);
inv M7_CSL0_CL2_LB1_Mux2_0(in265, M7_CSL0_CL2_LB1_Not_ContIn);
and2 M7_CSL0_CL2_LB1_Mux2_1(NotContLogic3_0_2, M7_CSL0_CL2_LB1_Not_ContIn, M7_CSL0_CL2_LB1_line1);
and2 M7_CSL0_CL2_LB1_Mux2_2(NotContLogic3_0_3, in265, M7_CSL0_CL2_LB1_line2);
or2 M7_CSL0_CL2_LB1_Mux2_3(M7_CSL0_CL2_LB1_line1, M7_CSL0_CL2_LB1_line2, M7_CSL0_CL2_line1);
or2 M7_CSL0_CL2_LB2(in400, M7_CSL0_CL2_line0, M7_CSL0_CL2_line2);
nand2 M7_CSL0_CL2_LB3(in400, M7_CSL0_CL2_line1, M7_CSL0_CL2_line3);
and2 M7_CSL0_CL2_LB4(M7_CSL0_CL2_line2, M7_CSL0_CL2_line3, LogicYbus_2);
inv M7_CSL0_CL3_LB0_Mux2_0(in257, M7_CSL0_CL3_LB0_Not_ContIn);
and2 M7_CSL0_CL3_LB0_Mux2_1(NotContLogic3_0_0, M7_CSL0_CL3_LB0_Not_ContIn, M7_CSL0_CL3_LB0_line1);
and2 M7_CSL0_CL3_LB0_Mux2_2(NotContLogic3_0_1, in257, M7_CSL0_CL3_LB0_line2);
or2 M7_CSL0_CL3_LB0_Mux2_3(M7_CSL0_CL3_LB0_line1, M7_CSL0_CL3_LB0_line2, M7_CSL0_CL3_line0);
inv M7_CSL0_CL3_LB1_Mux2_0(in257, M7_CSL0_CL3_LB1_Not_ContIn);
and2 M7_CSL0_CL3_LB1_Mux2_1(NotContLogic3_0_2, M7_CSL0_CL3_LB1_Not_ContIn, M7_CSL0_CL3_LB1_line1);
and2 M7_CSL0_CL3_LB1_Mux2_2(NotContLogic3_0_3, in257, M7_CSL0_CL3_LB1_line2);
or2 M7_CSL0_CL3_LB1_Mux2_3(M7_CSL0_CL3_LB1_line1, M7_CSL0_CL3_LB1_line2, M7_CSL0_CL3_line1);
or2 M7_CSL0_CL3_LB2(in389, M7_CSL0_CL3_line0, M7_CSL0_CL3_line2);
nand2 M7_CSL0_CL3_LB3(in389, M7_CSL0_CL3_line1, M7_CSL0_CL3_line3);
and2 M7_CSL0_CL3_LB4(M7_CSL0_CL3_line2, M7_CSL0_CL3_line3, LogicYbus_3);
inv M7_CSL0_CL4_LB0_Mux2_0(in234, M7_CSL0_CL4_LB0_Not_ContIn);
and2 M7_CSL0_CL4_LB0_Mux2_1(NotContLogic3_0_0, M7_CSL0_CL4_LB0_Not_ContIn, M7_CSL0_CL4_LB0_line1);
and2 M7_CSL0_CL4_LB0_Mux2_2(NotContLogic3_0_1, in234, M7_CSL0_CL4_LB0_line2);
or2 M7_CSL0_CL4_LB0_Mux2_3(M7_CSL0_CL4_LB0_line1, M7_CSL0_CL4_LB0_line2, M7_CSL0_CL4_line0);
inv M7_CSL0_CL4_LB1_Mux2_0(in234, M7_CSL0_CL4_LB1_Not_ContIn);
and2 M7_CSL0_CL4_LB1_Mux2_1(NotContLogic3_0_2, M7_CSL0_CL4_LB1_Not_ContIn, M7_CSL0_CL4_LB1_line1);
and2 M7_CSL0_CL4_LB1_Mux2_2(NotContLogic3_0_3, in234, M7_CSL0_CL4_LB1_line2);
or2 M7_CSL0_CL4_LB1_Mux2_3(M7_CSL0_CL4_LB1_line1, M7_CSL0_CL4_LB1_line2, M7_CSL0_CL4_line1);
or2 M7_CSL0_CL4_LB2(in435, M7_CSL0_CL4_line0, M7_CSL0_CL4_line2);
nand2 M7_CSL0_CL4_LB3(in435, M7_CSL0_CL4_line1, M7_CSL0_CL4_line3);
and2 M7_CSL0_CL4_LB4(M7_CSL0_CL4_line2, M7_CSL0_CL4_line3, LogicYbus_4);
inv M7_CSL0_CL5_LB0_Mux2_0(in226, M7_CSL0_CL5_LB0_Not_ContIn);
and2 M7_CSL0_CL5_LB0_Mux2_1(NotContLogic3_0_0, M7_CSL0_CL5_LB0_Not_ContIn, M7_CSL0_CL5_LB0_line1);
and2 M7_CSL0_CL5_LB0_Mux2_2(NotContLogic3_0_1, in226, M7_CSL0_CL5_LB0_line2);
or2 M7_CSL0_CL5_LB0_Mux2_3(M7_CSL0_CL5_LB0_line1, M7_CSL0_CL5_LB0_line2, M7_CSL0_CL5_line0);
inv M7_CSL0_CL5_LB1_Mux2_0(in226, M7_CSL0_CL5_LB1_Not_ContIn);
and2 M7_CSL0_CL5_LB1_Mux2_1(NotContLogic3_0_2, M7_CSL0_CL5_LB1_Not_ContIn, M7_CSL0_CL5_LB1_line1);
and2 M7_CSL0_CL5_LB1_Mux2_2(NotContLogic3_0_3, in226, M7_CSL0_CL5_LB1_line2);
or2 M7_CSL0_CL5_LB1_Mux2_3(M7_CSL0_CL5_LB1_line1, M7_CSL0_CL5_LB1_line2, M7_CSL0_CL5_line1);
or2 M7_CSL0_CL5_LB2(in422, M7_CSL0_CL5_line0, M7_CSL0_CL5_line2);
nand2 M7_CSL0_CL5_LB3(in422, M7_CSL0_CL5_line1, M7_CSL0_CL5_line3);
and2 M7_CSL0_CL5_LB4(M7_CSL0_CL5_line2, M7_CSL0_CL5_line3, LogicYbus_5);
inv M7_CSL0_CL6_LB0_Mux2_0(in218, M7_CSL0_CL6_LB0_Not_ContIn);
and2 M7_CSL0_CL6_LB0_Mux2_1(NotContLogic3_0_0, M7_CSL0_CL6_LB0_Not_ContIn, M7_CSL0_CL6_LB0_line1);
and2 M7_CSL0_CL6_LB0_Mux2_2(NotContLogic3_0_1, in218, M7_CSL0_CL6_LB0_line2);
or2 M7_CSL0_CL6_LB0_Mux2_3(M7_CSL0_CL6_LB0_line1, M7_CSL0_CL6_LB0_line2, M7_CSL0_CL6_line0);
inv M7_CSL0_CL6_LB1_Mux2_0(in218, M7_CSL0_CL6_LB1_Not_ContIn);
and2 M7_CSL0_CL6_LB1_Mux2_1(NotContLogic3_0_2, M7_CSL0_CL6_LB1_Not_ContIn, M7_CSL0_CL6_LB1_line1);
and2 M7_CSL0_CL6_LB1_Mux2_2(NotContLogic3_0_3, in218, M7_CSL0_CL6_LB1_line2);
or2 M7_CSL0_CL6_LB1_Mux2_3(M7_CSL0_CL6_LB1_line1, M7_CSL0_CL6_LB1_line2, M7_CSL0_CL6_line1);
or2 M7_CSL0_CL6_LB2(in468, M7_CSL0_CL6_line0, M7_CSL0_CL6_line2);
nand2 M7_CSL0_CL6_LB3(in468, M7_CSL0_CL6_line1, M7_CSL0_CL6_line3);
and2 M7_CSL0_CL6_LB4(M7_CSL0_CL6_line2, M7_CSL0_CL6_line3, LogicYbus_6);
inv M7_CSL0_CL7_LB0_Mux2_0(in210, M7_CSL0_CL7_LB0_Not_ContIn);
and2 M7_CSL0_CL7_LB0_Mux2_1(NotContLogic3_0_0, M7_CSL0_CL7_LB0_Not_ContIn, M7_CSL0_CL7_LB0_line1);
and2 M7_CSL0_CL7_LB0_Mux2_2(NotContLogic3_0_1, in210, M7_CSL0_CL7_LB0_line2);
or2 M7_CSL0_CL7_LB0_Mux2_3(M7_CSL0_CL7_LB0_line1, M7_CSL0_CL7_LB0_line2, M7_CSL0_CL7_line0);
inv M7_CSL0_CL7_LB1_Mux2_0(in210, M7_CSL0_CL7_LB1_Not_ContIn);
and2 M7_CSL0_CL7_LB1_Mux2_1(NotContLogic3_0_2, M7_CSL0_CL7_LB1_Not_ContIn, M7_CSL0_CL7_LB1_line1);
and2 M7_CSL0_CL7_LB1_Mux2_2(NotContLogic3_0_3, in210, M7_CSL0_CL7_LB1_line2);
or2 M7_CSL0_CL7_LB1_Mux2_3(M7_CSL0_CL7_LB1_line1, M7_CSL0_CL7_LB1_line2, M7_CSL0_CL7_line1);
or2 M7_CSL0_CL7_LB2(in457, M7_CSL0_CL7_line0, M7_CSL0_CL7_line2);
nand2 M7_CSL0_CL7_LB3(in457, M7_CSL0_CL7_line1, M7_CSL0_CL7_line3);
and2 M7_CSL0_CL7_LB4(M7_CSL0_CL7_line2, M7_CSL0_CL7_line3, LogicYbus_7);
inv M7_CSL0_CL8_LB0_Mux2_0(in206, M7_CSL0_CL8_LB0_Not_ContIn);
and2 M7_CSL0_CL8_LB0_Mux2_1(in254, M7_CSL0_CL8_LB0_Not_ContIn, M7_CSL0_CL8_LB0_line1);
and2 M7_CSL0_CL8_LB0_Mux2_2(in242, in206, M7_CSL0_CL8_LB0_line2);
or2 M7_CSL0_CL8_LB0_Mux2_3(M7_CSL0_CL8_LB0_line1, M7_CSL0_CL8_LB0_line2, M7_CSL0_CL8_line0);
inv M7_CSL0_CL8_LB1_Mux2_0(in206, M7_CSL0_CL8_LB1_Not_ContIn);
and2 M7_CSL0_CL8_LB1_Mux2_1(in251, M7_CSL0_CL8_LB1_Not_ContIn, M7_CSL0_CL8_LB1_line1);
and2 M7_CSL0_CL8_LB1_Mux2_2(in248, in206, M7_CSL0_CL8_LB1_line2);
or2 M7_CSL0_CL8_LB1_Mux2_3(M7_CSL0_CL8_LB1_line1, M7_CSL0_CL8_LB1_line2, M7_CSL0_CL8_line1);
or2 M7_CSL0_CL8_LB2(in446, M7_CSL0_CL8_line0, M7_CSL0_CL8_line2);
nand2 M7_CSL0_CL8_LB3(in446, M7_CSL0_CL8_line1, M7_CSL0_CL8_line3);
and2 M7_CSL0_CL8_LB4(M7_CSL0_CL8_line2, M7_CSL0_CL8_line3, LogicYbus_8);
and2 M7_CSL1_Add0_GP9_0(Ybus_0, in374, M7_CSL1_Genbus_0);
and2 M7_CSL1_Add0_GP9_1(Ybus_1, in411, M7_CSL1_Genbus_1);
and2 M7_CSL1_Add0_GP9_2(Ybus_2, in400, M7_CSL1_Genbus_2);
and2 M7_CSL1_Add0_GP9_3(Ybus_3, in389, M7_CSL1_Genbus_3);
and2 M7_CSL1_Add0_GP9_4(Ybus_4, in435, M7_CSL1_Genbus_4);
and2 M7_CSL1_Add0_GP9_5(Ybus_5, in422, M7_CSL1_Genbus_5);
and2 M7_CSL1_Add0_GP9_6(Ybus_6, in468, M7_CSL1_Genbus_6);
and2 M7_CSL1_Add0_GP9_7(Ybus_7, in457, M7_CSL1_Genbus_7);
and2 M7_CSL1_Add0_GP9_8(Ybus_8, in446, M7_CSL1_Genbus_8);
inv M7_CSL1_Add0_GP9_9_Xo0(Ybus_0, M7_CSL1_Add0_GP9_9_NotA);
inv M7_CSL1_Add0_GP9_9_Xo1(in374, M7_CSL1_Add0_GP9_9_NotB);
nand2 M7_CSL1_Add0_GP9_9_Xo2(M7_CSL1_Add0_GP9_9_NotA, in374, M7_CSL1_Add0_GP9_9_line2);
nand2 M7_CSL1_Add0_GP9_9_Xo3(M7_CSL1_Add0_GP9_9_NotB, Ybus_0, M7_CSL1_Add0_GP9_9_line3);
nand2 M7_CSL1_Add0_GP9_9_Xo4(M7_CSL1_Add0_GP9_9_line2, M7_CSL1_Add0_GP9_9_line3, M7_CSL1_Propbus_0);
inv M7_CSL1_Add0_GP9_10_Xo0(Ybus_1, M7_CSL1_Add0_GP9_10_NotA);
inv M7_CSL1_Add0_GP9_10_Xo1(in411, M7_CSL1_Add0_GP9_10_NotB);
nand2 M7_CSL1_Add0_GP9_10_Xo2(M7_CSL1_Add0_GP9_10_NotA, in411, M7_CSL1_Add0_GP9_10_line2);
nand2 M7_CSL1_Add0_GP9_10_Xo3(M7_CSL1_Add0_GP9_10_NotB, Ybus_1, M7_CSL1_Add0_GP9_10_line3);
nand2 M7_CSL1_Add0_GP9_10_Xo4(M7_CSL1_Add0_GP9_10_line2, M7_CSL1_Add0_GP9_10_line3, M7_CSL1_Propbus_1);
inv M7_CSL1_Add0_GP9_11_Xo0(Ybus_2, M7_CSL1_Add0_GP9_11_NotA);
inv M7_CSL1_Add0_GP9_11_Xo1(in400, M7_CSL1_Add0_GP9_11_NotB);
nand2 M7_CSL1_Add0_GP9_11_Xo2(M7_CSL1_Add0_GP9_11_NotA, in400, M7_CSL1_Add0_GP9_11_line2);
nand2 M7_CSL1_Add0_GP9_11_Xo3(M7_CSL1_Add0_GP9_11_NotB, Ybus_2, M7_CSL1_Add0_GP9_11_line3);
nand2 M7_CSL1_Add0_GP9_11_Xo4(M7_CSL1_Add0_GP9_11_line2, M7_CSL1_Add0_GP9_11_line3, M7_CSL1_Propbus_2);
inv M7_CSL1_Add0_GP9_12_Xo0(Ybus_3, M7_CSL1_Add0_GP9_12_NotA);
inv M7_CSL1_Add0_GP9_12_Xo1(in389, M7_CSL1_Add0_GP9_12_NotB);
nand2 M7_CSL1_Add0_GP9_12_Xo2(M7_CSL1_Add0_GP9_12_NotA, in389, M7_CSL1_Add0_GP9_12_line2);
nand2 M7_CSL1_Add0_GP9_12_Xo3(M7_CSL1_Add0_GP9_12_NotB, Ybus_3, M7_CSL1_Add0_GP9_12_line3);
nand2 M7_CSL1_Add0_GP9_12_Xo4(M7_CSL1_Add0_GP9_12_line2, M7_CSL1_Add0_GP9_12_line3, M7_CSL1_Propbus_3);
inv M7_CSL1_Add0_GP9_13_Xo0(Ybus_4, M7_CSL1_Add0_GP9_13_NotA);
inv M7_CSL1_Add0_GP9_13_Xo1(in435, M7_CSL1_Add0_GP9_13_NotB);
nand2 M7_CSL1_Add0_GP9_13_Xo2(M7_CSL1_Add0_GP9_13_NotA, in435, M7_CSL1_Add0_GP9_13_line2);
nand2 M7_CSL1_Add0_GP9_13_Xo3(M7_CSL1_Add0_GP9_13_NotB, Ybus_4, M7_CSL1_Add0_GP9_13_line3);
nand2 M7_CSL1_Add0_GP9_13_Xo4(M7_CSL1_Add0_GP9_13_line2, M7_CSL1_Add0_GP9_13_line3, M7_CSL1_Propbus_4);
inv M7_CSL1_Add0_GP9_14_Xo0(Ybus_5, M7_CSL1_Add0_GP9_14_NotA);
inv M7_CSL1_Add0_GP9_14_Xo1(in422, M7_CSL1_Add0_GP9_14_NotB);
nand2 M7_CSL1_Add0_GP9_14_Xo2(M7_CSL1_Add0_GP9_14_NotA, in422, M7_CSL1_Add0_GP9_14_line2);
nand2 M7_CSL1_Add0_GP9_14_Xo3(M7_CSL1_Add0_GP9_14_NotB, Ybus_5, M7_CSL1_Add0_GP9_14_line3);
nand2 M7_CSL1_Add0_GP9_14_Xo4(M7_CSL1_Add0_GP9_14_line2, M7_CSL1_Add0_GP9_14_line3, M7_CSL1_Propbus_5);
inv M7_CSL1_Add0_GP9_15_Xo0(Ybus_6, M7_CSL1_Add0_GP9_15_NotA);
inv M7_CSL1_Add0_GP9_15_Xo1(in468, M7_CSL1_Add0_GP9_15_NotB);
nand2 M7_CSL1_Add0_GP9_15_Xo2(M7_CSL1_Add0_GP9_15_NotA, in468, M7_CSL1_Add0_GP9_15_line2);
nand2 M7_CSL1_Add0_GP9_15_Xo3(M7_CSL1_Add0_GP9_15_NotB, Ybus_6, M7_CSL1_Add0_GP9_15_line3);
nand2 M7_CSL1_Add0_GP9_15_Xo4(M7_CSL1_Add0_GP9_15_line2, M7_CSL1_Add0_GP9_15_line3, M7_CSL1_Propbus_6);
inv M7_CSL1_Add0_GP9_16_Xo0(Ybus_7, M7_CSL1_Add0_GP9_16_NotA);
inv M7_CSL1_Add0_GP9_16_Xo1(in457, M7_CSL1_Add0_GP9_16_NotB);
nand2 M7_CSL1_Add0_GP9_16_Xo2(M7_CSL1_Add0_GP9_16_NotA, in457, M7_CSL1_Add0_GP9_16_line2);
nand2 M7_CSL1_Add0_GP9_16_Xo3(M7_CSL1_Add0_GP9_16_NotB, Ybus_7, M7_CSL1_Add0_GP9_16_line3);
nand2 M7_CSL1_Add0_GP9_16_Xo4(M7_CSL1_Add0_GP9_16_line2, M7_CSL1_Add0_GP9_16_line3, M7_CSL1_Propbus_7);
inv M7_CSL1_Add0_GP9_17_Xo0(Ybus_8, M7_CSL1_Add0_GP9_17_NotA);
inv M7_CSL1_Add0_GP9_17_Xo1(in446, M7_CSL1_Add0_GP9_17_NotB);
nand2 M7_CSL1_Add0_GP9_17_Xo2(M7_CSL1_Add0_GP9_17_NotA, in446, M7_CSL1_Add0_GP9_17_line2);
nand2 M7_CSL1_Add0_GP9_17_Xo3(M7_CSL1_Add0_GP9_17_NotB, Ybus_8, M7_CSL1_Add0_GP9_17_line3);
nand2 M7_CSL1_Add0_GP9_17_Xo4(M7_CSL1_Add0_GP9_17_line2, M7_CSL1_Add0_GP9_17_line3, M7_CSL1_Propbus_8);
and2 M7_CSL1_Add1_CB0_Ao2_0(M7_CSL1_Propbus_0, in4, M7_CSL1_Add1_CB0_line0);
or2 M7_CSL1_Add1_CB0_Ao2_1(M7_CSL1_Genbus_0, M7_CSL1_Add1_CB0_line0, M7_CSL1_Carry_0);
and2 M7_CSL1_Add1_CB1_Ao3a_0(M7_CSL1_Propbus_1, M7_CSL1_Genbus_0, M7_CSL1_Add1_CB1_line0);
and3 M7_CSL1_Add1_CB1_Ao3a_1(M7_CSL1_Propbus_1, M7_CSL1_Propbus_0, in4, M7_CSL1_Add1_CB1_line1);
or3 M7_CSL1_Add1_CB1_Ao3a_2(M7_CSL1_Genbus_1, M7_CSL1_Add1_CB1_line0, M7_CSL1_Add1_CB1_line1, M7_CSL1_Carry_1);
and2 M7_CSL1_Add1_CB2_Ao4a_0(M7_CSL1_Propbus_2, M7_CSL1_Genbus_1, M7_CSL1_Add1_CB2_line0);
and3 M7_CSL1_Add1_CB2_Ao4a_1(M7_CSL1_Propbus_2, M7_CSL1_Propbus_1, M7_CSL1_Genbus_0, M7_CSL1_Add1_CB2_line1);
and4 M7_CSL1_Add1_CB2_Ao4a_2(M7_CSL1_Propbus_2, M7_CSL1_Propbus_1, M7_CSL1_Propbus_0, in4, M7_CSL1_Add1_CB2_line2);
or4 M7_CSL1_Add1_CB2_Ao4a_3(M7_CSL1_Genbus_2, M7_CSL1_Add1_CB2_line0, M7_CSL1_Add1_CB2_line1, M7_CSL1_Add1_CB2_line2, M7_CSL1_Carry_2);
and2 M7_CSL1_Add1_CB3_Ao5a_0(M7_CSL1_Propbus_3, M7_CSL1_Genbus_2, M7_CSL1_Add1_CB3_line0);
and3 M7_CSL1_Add1_CB3_Ao5a_1(M7_CSL1_Propbus_3, M7_CSL1_Propbus_2, M7_CSL1_Genbus_1, M7_CSL1_Add1_CB3_line1);
and4 M7_CSL1_Add1_CB3_Ao5a_2(M7_CSL1_Propbus_3, M7_CSL1_Propbus_2, M7_CSL1_Propbus_1, M7_CSL1_Genbus_0, M7_CSL1_Add1_CB3_line2);
and5 M7_CSL1_Add1_CB3_Ao5a_3(M7_CSL1_Propbus_3, M7_CSL1_Propbus_2, M7_CSL1_Propbus_1, M7_CSL1_Propbus_0, in4, M7_CSL1_Add1_CB3_line3);
or5 M7_CSL1_Add1_CB3_Ao5a_4(M7_CSL1_Genbus_3, M7_CSL1_Add1_CB3_line0, M7_CSL1_Add1_CB3_line1, M7_CSL1_Add1_CB3_line2, M7_CSL1_Add1_CB3_line3, M7_CSL1_Carry_3);
and2 M7_CSL1_Add1_CB4_Ao5a_0(M7_CSL1_Propbus_4, M7_CSL1_Genbus_3, M7_CSL1_Add1_CB4_line0);
and3 M7_CSL1_Add1_CB4_Ao5a_1(M7_CSL1_Propbus_4, M7_CSL1_Propbus_3, M7_CSL1_Genbus_2, M7_CSL1_Add1_CB4_line1);
and4 M7_CSL1_Add1_CB4_Ao5a_2(M7_CSL1_Propbus_4, M7_CSL1_Propbus_3, M7_CSL1_Propbus_2, M7_CSL1_Genbus_1, M7_CSL1_Add1_CB4_line2);
and5 M7_CSL1_Add1_CB4_Ao5a_3(M7_CSL1_Propbus_4, M7_CSL1_Propbus_3, M7_CSL1_Propbus_2, M7_CSL1_Propbus_1, M7_CSL1_Genbus_0, M7_CSL1_Add1_CB4_line3);
or5 M7_CSL1_Add1_CB4_Ao5a_4(M7_CSL1_Genbus_4, M7_CSL1_Add1_CB4_line0, M7_CSL1_Add1_CB4_line1, M7_CSL1_Add1_CB4_line2, M7_CSL1_Add1_CB4_line3, M7_CSL1_Add1_LocalC0_4);
and5 M7_CSL1_Add1_CB5(M7_CSL1_Propbus_0, M7_CSL1_Propbus_1, M7_CSL1_Propbus_2, M7_CSL1_Propbus_3, M7_CSL1_Propbus_4, M7_CSL1_Add1_Prop4_0);
and2 M7_CSL1_Add1_CB6(in4, M7_CSL1_Add1_Prop4_0, M7_CSL1_Add1_PropCin);
or2 M7_CSL1_Add1_CB7(M7_CSL1_Add1_LocalC0_4, M7_CSL1_Add1_PropCin, M7_CSL1_Carry_4);
and2 M7_CSL1_Add1_CB8_Ao5a_0(M7_CSL1_Propbus_8, M7_CSL1_Genbus_7, M7_CSL1_Add1_CB8_line0);
and3 M7_CSL1_Add1_CB8_Ao5a_1(M7_CSL1_Propbus_8, M7_CSL1_Propbus_7, M7_CSL1_Genbus_6, M7_CSL1_Add1_CB8_line1);
and4 M7_CSL1_Add1_CB8_Ao5a_2(M7_CSL1_Propbus_8, M7_CSL1_Propbus_7, M7_CSL1_Propbus_6, M7_CSL1_Genbus_5, M7_CSL1_Add1_CB8_line2);
and5 M7_CSL1_Add1_CB8_Ao5a_3(M7_CSL1_Propbus_8, M7_CSL1_Propbus_7, M7_CSL1_Propbus_6, M7_CSL1_Propbus_5, M7_CSL1_Add1_LocalC0_4, M7_CSL1_Add1_CB8_line3);
or5 M7_CSL1_Add1_CB8_Ao5a_4(M7_CSL1_Genbus_8, M7_CSL1_Add1_CB8_line0, M7_CSL1_Add1_CB8_line1, M7_CSL1_Add1_CB8_line2, M7_CSL1_Add1_CB8_line3, out591);
and4 M7_CSL1_Add1_CB9(M7_CSL1_Propbus_5, M7_CSL1_Propbus_6, M7_CSL1_Propbus_7, M7_CSL1_Propbus_8, M7_CSL1_Add1_Prop8_5);
and2 M7_CSL1_Add1_CB10(M7_CSL1_Add1_Prop4_0, M7_CSL1_Add1_Prop8_5, out588);
or2 M7_CSL1_Add2_GLC4_0(M7_CSL1_Genbus_5, M7_CSL1_Propbus_5, M7_CSL1_LocalHC1_0);
and2 M7_CSL1_Add2_GLC4_1_Ao2_0(M7_CSL1_Propbus_6, M7_CSL1_Genbus_5, M7_CSL1_Add2_GLC4_1_line0);
or2 M7_CSL1_Add2_GLC4_1_Ao2_1(M7_CSL1_Genbus_6, M7_CSL1_Add2_GLC4_1_line0, M7_CSL1_LocalHC0_1);
and2 M7_CSL1_Add2_GLC4_2_Ao3a_0(M7_CSL1_Propbus_6, M7_CSL1_Genbus_5, M7_CSL1_Add2_GLC4_2_line0);
and2 M7_CSL1_Add2_GLC4_2_Ao3a_1(M7_CSL1_Propbus_6, M7_CSL1_Propbus_5, M7_CSL1_Add2_GLC4_2_line1);
or3 M7_CSL1_Add2_GLC4_2_Ao3a_2(M7_CSL1_Genbus_6, M7_CSL1_Add2_GLC4_2_line0, M7_CSL1_Add2_GLC4_2_line1, M7_CSL1_LocalHC1_1);
and2 M7_CSL1_Add2_GLC4_3_Ao3a_0(M7_CSL1_Propbus_7, M7_CSL1_Genbus_6, M7_CSL1_Add2_GLC4_3_line0);
and3 M7_CSL1_Add2_GLC4_3_Ao3a_1(M7_CSL1_Propbus_7, M7_CSL1_Propbus_6, M7_CSL1_Genbus_5, M7_CSL1_Add2_GLC4_3_line1);
or3 M7_CSL1_Add2_GLC4_3_Ao3a_2(M7_CSL1_Genbus_7, M7_CSL1_Add2_GLC4_3_line0, M7_CSL1_Add2_GLC4_3_line1, M7_CSL1_LocalHC0_2);
and2 M7_CSL1_Add2_GLC4_4_Ao4a_0(M7_CSL1_Propbus_7, M7_CSL1_Genbus_6, M7_CSL1_Add2_GLC4_4_line0);
and3 M7_CSL1_Add2_GLC4_4_Ao4a_1(M7_CSL1_Propbus_7, M7_CSL1_Propbus_6, M7_CSL1_Genbus_5, M7_CSL1_Add2_GLC4_4_line1);
and3 M7_CSL1_Add2_GLC4_4_Ao4a_2(M7_CSL1_Propbus_7, M7_CSL1_Propbus_6, M7_CSL1_Propbus_5, M7_CSL1_Add2_GLC4_4_line2);
or4 M7_CSL1_Add2_GLC4_4_Ao4a_3(M7_CSL1_Genbus_7, M7_CSL1_Add2_GLC4_4_line0, M7_CSL1_Add2_GLC4_4_line1, M7_CSL1_Add2_GLC4_4_line2, M7_CSL1_LocalHC1_2);
inv M7_CSL1_Add3_X2a6_0_Xo0(M7_CSL1_Propbus_0, M7_CSL1_Add3_X2a6_0_NotA);
inv M7_CSL1_Add3_X2a6_0_Xo1(in4, M7_CSL1_Add3_X2a6_0_NotB);
nand2 M7_CSL1_Add3_X2a6_0_Xo2(M7_CSL1_Add3_X2a6_0_NotA, in4, M7_CSL1_Add3_X2a6_0_line2);
nand2 M7_CSL1_Add3_X2a6_0_Xo3(M7_CSL1_Add3_X2a6_0_NotB, M7_CSL1_Propbus_0, M7_CSL1_Add3_X2a6_0_line3);
nand2 M7_CSL1_Add3_X2a6_0_Xo4(M7_CSL1_Add3_X2a6_0_line2, M7_CSL1_Add3_X2a6_0_line3, SumYbus_0);
inv M7_CSL1_Add3_X2a6_1_Xo0(M7_CSL1_Propbus_1, M7_CSL1_Add3_X2a6_1_NotA);
inv M7_CSL1_Add3_X2a6_1_Xo1(M7_CSL1_Carry_0, M7_CSL1_Add3_X2a6_1_NotB);
nand2 M7_CSL1_Add3_X2a6_1_Xo2(M7_CSL1_Add3_X2a6_1_NotA, M7_CSL1_Carry_0, M7_CSL1_Add3_X2a6_1_line2);
nand2 M7_CSL1_Add3_X2a6_1_Xo3(M7_CSL1_Add3_X2a6_1_NotB, M7_CSL1_Propbus_1, M7_CSL1_Add3_X2a6_1_line3);
nand2 M7_CSL1_Add3_X2a6_1_Xo4(M7_CSL1_Add3_X2a6_1_line2, M7_CSL1_Add3_X2a6_1_line3, SumYbus_1);
inv M7_CSL1_Add3_X2a6_2_Xo0(M7_CSL1_Propbus_2, M7_CSL1_Add3_X2a6_2_NotA);
inv M7_CSL1_Add3_X2a6_2_Xo1(M7_CSL1_Carry_1, M7_CSL1_Add3_X2a6_2_NotB);
nand2 M7_CSL1_Add3_X2a6_2_Xo2(M7_CSL1_Add3_X2a6_2_NotA, M7_CSL1_Carry_1, M7_CSL1_Add3_X2a6_2_line2);
nand2 M7_CSL1_Add3_X2a6_2_Xo3(M7_CSL1_Add3_X2a6_2_NotB, M7_CSL1_Propbus_2, M7_CSL1_Add3_X2a6_2_line3);
nand2 M7_CSL1_Add3_X2a6_2_Xo4(M7_CSL1_Add3_X2a6_2_line2, M7_CSL1_Add3_X2a6_2_line3, SumYbus_2);
inv M7_CSL1_Add3_X2a6_3_Xo0(M7_CSL1_Propbus_3, M7_CSL1_Add3_X2a6_3_NotA);
inv M7_CSL1_Add3_X2a6_3_Xo1(M7_CSL1_Carry_2, M7_CSL1_Add3_X2a6_3_NotB);
nand2 M7_CSL1_Add3_X2a6_3_Xo2(M7_CSL1_Add3_X2a6_3_NotA, M7_CSL1_Carry_2, M7_CSL1_Add3_X2a6_3_line2);
nand2 M7_CSL1_Add3_X2a6_3_Xo3(M7_CSL1_Add3_X2a6_3_NotB, M7_CSL1_Propbus_3, M7_CSL1_Add3_X2a6_3_line3);
nand2 M7_CSL1_Add3_X2a6_3_Xo4(M7_CSL1_Add3_X2a6_3_line2, M7_CSL1_Add3_X2a6_3_line3, SumYbus_3);
inv M7_CSL1_Add3_X2a6_4_Xo0(M7_CSL1_Propbus_4, M7_CSL1_Add3_X2a6_4_NotA);
inv M7_CSL1_Add3_X2a6_4_Xo1(M7_CSL1_Carry_3, M7_CSL1_Add3_X2a6_4_NotB);
nand2 M7_CSL1_Add3_X2a6_4_Xo2(M7_CSL1_Add3_X2a6_4_NotA, M7_CSL1_Carry_3, M7_CSL1_Add3_X2a6_4_line2);
nand2 M7_CSL1_Add3_X2a6_4_Xo3(M7_CSL1_Add3_X2a6_4_NotB, M7_CSL1_Propbus_4, M7_CSL1_Add3_X2a6_4_line3);
nand2 M7_CSL1_Add3_X2a6_4_Xo4(M7_CSL1_Add3_X2a6_4_line2, M7_CSL1_Add3_X2a6_4_line3, SumYbus_4);
inv M7_CSL1_Add3_X2a6_5_Xo0(M7_CSL1_Propbus_5, M7_CSL1_Add3_X2a6_5_NotA);
inv M7_CSL1_Add3_X2a6_5_Xo1(M7_CSL1_Carry_4, M7_CSL1_Add3_X2a6_5_NotB);
nand2 M7_CSL1_Add3_X2a6_5_Xo2(M7_CSL1_Add3_X2a6_5_NotA, M7_CSL1_Carry_4, M7_CSL1_Add3_X2a6_5_line2);
nand2 M7_CSL1_Add3_X2a6_5_Xo3(M7_CSL1_Add3_X2a6_5_NotB, M7_CSL1_Propbus_5, M7_CSL1_Add3_X2a6_5_line3);
nand2 M7_CSL1_Add3_X2a6_5_Xo4(M7_CSL1_Add3_X2a6_5_line2, M7_CSL1_Add3_X2a6_5_line3, SumYbus_5);
inv M7_CSL1_Add4_X2a6_0_Xo0(M7_CSL1_Propbus_6, M7_CSL1_Add4_X2a6_0_NotA);
inv M7_CSL1_Add4_X2a6_0_Xo1(M7_CSL1_Genbus_5, M7_CSL1_Add4_X2a6_0_NotB);
nand2 M7_CSL1_Add4_X2a6_0_Xo2(M7_CSL1_Add4_X2a6_0_NotA, M7_CSL1_Genbus_5, M7_CSL1_Add4_X2a6_0_line2);
nand2 M7_CSL1_Add4_X2a6_0_Xo3(M7_CSL1_Add4_X2a6_0_NotB, M7_CSL1_Propbus_6, M7_CSL1_Add4_X2a6_0_line3);
nand2 M7_CSL1_Add4_X2a6_0_Xo4(M7_CSL1_Add4_X2a6_0_line2, M7_CSL1_Add4_X2a6_0_line3, M7_CSL1_SumH01bus_0);
inv M7_CSL1_Add4_X2a6_1_Xo0(M7_CSL1_Propbus_7, M7_CSL1_Add4_X2a6_1_NotA);
inv M7_CSL1_Add4_X2a6_1_Xo1(M7_CSL1_LocalHC0_1, M7_CSL1_Add4_X2a6_1_NotB);
nand2 M7_CSL1_Add4_X2a6_1_Xo2(M7_CSL1_Add4_X2a6_1_NotA, M7_CSL1_LocalHC0_1, M7_CSL1_Add4_X2a6_1_line2);
nand2 M7_CSL1_Add4_X2a6_1_Xo3(M7_CSL1_Add4_X2a6_1_NotB, M7_CSL1_Propbus_7, M7_CSL1_Add4_X2a6_1_line3);
nand2 M7_CSL1_Add4_X2a6_1_Xo4(M7_CSL1_Add4_X2a6_1_line2, M7_CSL1_Add4_X2a6_1_line3, M7_CSL1_SumH01bus_1);
inv M7_CSL1_Add4_X2a6_2_Xo0(M7_CSL1_Propbus_8, M7_CSL1_Add4_X2a6_2_NotA);
inv M7_CSL1_Add4_X2a6_2_Xo1(M7_CSL1_LocalHC0_2, M7_CSL1_Add4_X2a6_2_NotB);
nand2 M7_CSL1_Add4_X2a6_2_Xo2(M7_CSL1_Add4_X2a6_2_NotA, M7_CSL1_LocalHC0_2, M7_CSL1_Add4_X2a6_2_line2);
nand2 M7_CSL1_Add4_X2a6_2_Xo3(M7_CSL1_Add4_X2a6_2_NotB, M7_CSL1_Propbus_8, M7_CSL1_Add4_X2a6_2_line3);
nand2 M7_CSL1_Add4_X2a6_2_Xo4(M7_CSL1_Add4_X2a6_2_line2, M7_CSL1_Add4_X2a6_2_line3, M7_CSL1_SumH01bus_2);
inv M7_CSL1_Add4_X2a6_3_Xo0(M7_CSL1_Propbus_6, M7_CSL1_Add4_X2a6_3_NotA);
inv M7_CSL1_Add4_X2a6_3_Xo1(M7_CSL1_LocalHC1_0, M7_CSL1_Add4_X2a6_3_NotB);
nand2 M7_CSL1_Add4_X2a6_3_Xo2(M7_CSL1_Add4_X2a6_3_NotA, M7_CSL1_LocalHC1_0, M7_CSL1_Add4_X2a6_3_line2);
nand2 M7_CSL1_Add4_X2a6_3_Xo3(M7_CSL1_Add4_X2a6_3_NotB, M7_CSL1_Propbus_6, M7_CSL1_Add4_X2a6_3_line3);
nand2 M7_CSL1_Add4_X2a6_3_Xo4(M7_CSL1_Add4_X2a6_3_line2, M7_CSL1_Add4_X2a6_3_line3, M7_CSL1_SumH01bus_3);
inv M7_CSL1_Add4_X2a6_4_Xo0(M7_CSL1_Propbus_7, M7_CSL1_Add4_X2a6_4_NotA);
inv M7_CSL1_Add4_X2a6_4_Xo1(M7_CSL1_LocalHC1_1, M7_CSL1_Add4_X2a6_4_NotB);
nand2 M7_CSL1_Add4_X2a6_4_Xo2(M7_CSL1_Add4_X2a6_4_NotA, M7_CSL1_LocalHC1_1, M7_CSL1_Add4_X2a6_4_line2);
nand2 M7_CSL1_Add4_X2a6_4_Xo3(M7_CSL1_Add4_X2a6_4_NotB, M7_CSL1_Propbus_7, M7_CSL1_Add4_X2a6_4_line3);
nand2 M7_CSL1_Add4_X2a6_4_Xo4(M7_CSL1_Add4_X2a6_4_line2, M7_CSL1_Add4_X2a6_4_line3, M7_CSL1_SumH01bus_4);
inv M7_CSL1_Add4_X2a6_5_Xo0(M7_CSL1_Propbus_8, M7_CSL1_Add4_X2a6_5_NotA);
inv M7_CSL1_Add4_X2a6_5_Xo1(M7_CSL1_LocalHC1_2, M7_CSL1_Add4_X2a6_5_NotB);
nand2 M7_CSL1_Add4_X2a6_5_Xo2(M7_CSL1_Add4_X2a6_5_NotA, M7_CSL1_LocalHC1_2, M7_CSL1_Add4_X2a6_5_line2);
nand2 M7_CSL1_Add4_X2a6_5_Xo3(M7_CSL1_Add4_X2a6_5_NotB, M7_CSL1_Propbus_8, M7_CSL1_Add4_X2a6_5_line3);
nand2 M7_CSL1_Add4_X2a6_5_Xo4(M7_CSL1_Add4_X2a6_5_line2, M7_CSL1_Add4_X2a6_5_line3, M7_CSL1_SumH01bus_5);
inv M7_CSL1_Add5_Mux2_0(M7_CSL1_Carry_4, M7_CSL1_Add5_Not_ContIn);
and2 M7_CSL1_Add5_Mux2_1(M7_CSL1_SumH01bus_0, M7_CSL1_Add5_Not_ContIn, M7_CSL1_Add5_line1);
and2 M7_CSL1_Add5_Mux2_2(M7_CSL1_SumH01bus_3, M7_CSL1_Carry_4, M7_CSL1_Add5_line2);
or2 M7_CSL1_Add5_Mux2_3(M7_CSL1_Add5_line1, M7_CSL1_Add5_line2, SumYbus_6);
inv M7_CSL1_Add6_Mux2_0(M7_CSL1_Carry_4, M7_CSL1_Add6_Not_ContIn);
and2 M7_CSL1_Add6_Mux2_1(M7_CSL1_SumH01bus_1, M7_CSL1_Add6_Not_ContIn, M7_CSL1_Add6_line1);
and2 M7_CSL1_Add6_Mux2_2(M7_CSL1_SumH01bus_4, M7_CSL1_Carry_4, M7_CSL1_Add6_line2);
or2 M7_CSL1_Add6_Mux2_3(M7_CSL1_Add6_line1, M7_CSL1_Add6_line2, SumYbus_7);
inv M7_CSL1_Add7_Mux2_0(M7_CSL1_Carry_4, M7_CSL1_Add7_Not_ContIn);
and2 M7_CSL1_Add7_Mux2_1(M7_CSL1_SumH01bus_2, M7_CSL1_Add7_Not_ContIn, M7_CSL1_Add7_line1);
and2 M7_CSL1_Add7_Mux2_2(M7_CSL1_SumH01bus_5, M7_CSL1_Carry_4, M7_CSL1_Add7_line2);
or2 M7_CSL1_Add7_Mux2_3(M7_CSL1_Add7_line1, M7_CSL1_Add7_line2, SumYbus_8);
inv M7_CSL2_Mx9_0_Mx4_0_Mux4_0(in4092, M7_CSL2_Mx9_0_Mx4_0_Not_ContLo);
inv M7_CSL2_Mx9_0_Mx4_0_Mux4_1(in4091, M7_CSL2_Mx9_0_Mx4_0_Not_ContHi);
and3 M7_CSL2_Mx9_0_Mx4_0_Mux4_2(LogicYbus_0, M7_CSL2_Mx9_0_Mx4_0_Not_ContHi, M7_CSL2_Mx9_0_Mx4_0_Not_ContLo, M7_CSL2_Mx9_0_Mx4_0_line2);
and3 M7_CSL2_Mx9_0_Mx4_0_Mux4_3(in117, M7_CSL2_Mx9_0_Mx4_0_Not_ContHi, in4092, M7_CSL2_Mx9_0_Mx4_0_line3);
and3 M7_CSL2_Mx9_0_Mx4_0_Mux4_4(SumYbus_0, in4091, M7_CSL2_Mx9_0_Mx4_0_Not_ContLo, M7_CSL2_Mx9_0_Mx4_0_line4);
and3 M7_CSL2_Mx9_0_Mx4_0_Mux4_5(gnd, in4091, in4092, M7_CSL2_Mx9_0_Mx4_0_line5);
or4 M7_CSL2_Mx9_0_Mx4_0_Mux4_6(M7_CSL2_Mx9_0_Mx4_0_line2, M7_CSL2_Mx9_0_Mx4_0_line3, M7_CSL2_Mx9_0_Mx4_0_line4, M7_CSL2_Mx9_0_Mx4_0_line5, FYbus_0);
inv M7_CSL2_Mx9_0_Mx4_1_Mux4_0(in4092, M7_CSL2_Mx9_0_Mx4_1_Not_ContLo);
inv M7_CSL2_Mx9_0_Mx4_1_Mux4_1(in4091, M7_CSL2_Mx9_0_Mx4_1_Not_ContHi);
and3 M7_CSL2_Mx9_0_Mx4_1_Mux4_2(LogicYbus_1, M7_CSL2_Mx9_0_Mx4_1_Not_ContHi, M7_CSL2_Mx9_0_Mx4_1_Not_ContLo, M7_CSL2_Mx9_0_Mx4_1_line2);
and3 M7_CSL2_Mx9_0_Mx4_1_Mux4_3(in126, M7_CSL2_Mx9_0_Mx4_1_Not_ContHi, in4092, M7_CSL2_Mx9_0_Mx4_1_line3);
and3 M7_CSL2_Mx9_0_Mx4_1_Mux4_4(SumYbus_1, in4091, M7_CSL2_Mx9_0_Mx4_1_Not_ContLo, M7_CSL2_Mx9_0_Mx4_1_line4);
and3 M7_CSL2_Mx9_0_Mx4_1_Mux4_5(gnd, in4091, in4092, M7_CSL2_Mx9_0_Mx4_1_line5);
or4 M7_CSL2_Mx9_0_Mx4_1_Mux4_6(M7_CSL2_Mx9_0_Mx4_1_line2, M7_CSL2_Mx9_0_Mx4_1_line3, M7_CSL2_Mx9_0_Mx4_1_line4, M7_CSL2_Mx9_0_Mx4_1_line5, FYbus_1);
inv M7_CSL2_Mx9_0_Mx4_2_Mux4_0(in4092, M7_CSL2_Mx9_0_Mx4_2_Not_ContLo);
inv M7_CSL2_Mx9_0_Mx4_2_Mux4_1(in4091, M7_CSL2_Mx9_0_Mx4_2_Not_ContHi);
and3 M7_CSL2_Mx9_0_Mx4_2_Mux4_2(LogicYbus_2, M7_CSL2_Mx9_0_Mx4_2_Not_ContHi, M7_CSL2_Mx9_0_Mx4_2_Not_ContLo, M7_CSL2_Mx9_0_Mx4_2_line2);
and3 M7_CSL2_Mx9_0_Mx4_2_Mux4_3(in127, M7_CSL2_Mx9_0_Mx4_2_Not_ContHi, in4092, M7_CSL2_Mx9_0_Mx4_2_line3);
and3 M7_CSL2_Mx9_0_Mx4_2_Mux4_4(SumYbus_2, in4091, M7_CSL2_Mx9_0_Mx4_2_Not_ContLo, M7_CSL2_Mx9_0_Mx4_2_line4);
and3 M7_CSL2_Mx9_0_Mx4_2_Mux4_5(gnd, in4091, in4092, M7_CSL2_Mx9_0_Mx4_2_line5);
or4 M7_CSL2_Mx9_0_Mx4_2_Mux4_6(M7_CSL2_Mx9_0_Mx4_2_line2, M7_CSL2_Mx9_0_Mx4_2_line3, M7_CSL2_Mx9_0_Mx4_2_line4, M7_CSL2_Mx9_0_Mx4_2_line5, FYbus_2);
inv M7_CSL2_Mx9_0_Mx4_3_Mux4_0(in4092, M7_CSL2_Mx9_0_Mx4_3_Not_ContLo);
inv M7_CSL2_Mx9_0_Mx4_3_Mux4_1(in4091, M7_CSL2_Mx9_0_Mx4_3_Not_ContHi);
and3 M7_CSL2_Mx9_0_Mx4_3_Mux4_2(LogicYbus_3, M7_CSL2_Mx9_0_Mx4_3_Not_ContHi, M7_CSL2_Mx9_0_Mx4_3_Not_ContLo, M7_CSL2_Mx9_0_Mx4_3_line2);
and3 M7_CSL2_Mx9_0_Mx4_3_Mux4_3(in128, M7_CSL2_Mx9_0_Mx4_3_Not_ContHi, in4092, M7_CSL2_Mx9_0_Mx4_3_line3);
and3 M7_CSL2_Mx9_0_Mx4_3_Mux4_4(SumYbus_3, in4091, M7_CSL2_Mx9_0_Mx4_3_Not_ContLo, M7_CSL2_Mx9_0_Mx4_3_line4);
and3 M7_CSL2_Mx9_0_Mx4_3_Mux4_5(gnd, in4091, in4092, M7_CSL2_Mx9_0_Mx4_3_line5);
or4 M7_CSL2_Mx9_0_Mx4_3_Mux4_6(M7_CSL2_Mx9_0_Mx4_3_line2, M7_CSL2_Mx9_0_Mx4_3_line3, M7_CSL2_Mx9_0_Mx4_3_line4, M7_CSL2_Mx9_0_Mx4_3_line5, FYbus_3);
inv M7_CSL2_Mx9_1_Mx4_0_Mux4_0(in4092, M7_CSL2_Mx9_1_Mx4_0_Not_ContLo);
inv M7_CSL2_Mx9_1_Mx4_0_Mux4_1(in4091, M7_CSL2_Mx9_1_Mx4_0_Not_ContHi);
and3 M7_CSL2_Mx9_1_Mx4_0_Mux4_2(LogicYbus_4, M7_CSL2_Mx9_1_Mx4_0_Not_ContHi, M7_CSL2_Mx9_1_Mx4_0_Not_ContLo, M7_CSL2_Mx9_1_Mx4_0_line2);
and3 M7_CSL2_Mx9_1_Mx4_0_Mux4_3(in122, M7_CSL2_Mx9_1_Mx4_0_Not_ContHi, in4092, M7_CSL2_Mx9_1_Mx4_0_line3);
and3 M7_CSL2_Mx9_1_Mx4_0_Mux4_4(SumYbus_4, in4091, M7_CSL2_Mx9_1_Mx4_0_Not_ContLo, M7_CSL2_Mx9_1_Mx4_0_line4);
and3 M7_CSL2_Mx9_1_Mx4_0_Mux4_5(gnd, in4091, in4092, M7_CSL2_Mx9_1_Mx4_0_line5);
or4 M7_CSL2_Mx9_1_Mx4_0_Mux4_6(M7_CSL2_Mx9_1_Mx4_0_line2, M7_CSL2_Mx9_1_Mx4_0_line3, M7_CSL2_Mx9_1_Mx4_0_line4, M7_CSL2_Mx9_1_Mx4_0_line5, FYbus_4);
inv M7_CSL2_Mx9_1_Mx4_1_Mux4_0(in4092, M7_CSL2_Mx9_1_Mx4_1_Not_ContLo);
inv M7_CSL2_Mx9_1_Mx4_1_Mux4_1(in4091, M7_CSL2_Mx9_1_Mx4_1_Not_ContHi);
and3 M7_CSL2_Mx9_1_Mx4_1_Mux4_2(LogicYbus_5, M7_CSL2_Mx9_1_Mx4_1_Not_ContHi, M7_CSL2_Mx9_1_Mx4_1_Not_ContLo, M7_CSL2_Mx9_1_Mx4_1_line2);
and3 M7_CSL2_Mx9_1_Mx4_1_Mux4_3(in113, M7_CSL2_Mx9_1_Mx4_1_Not_ContHi, in4092, M7_CSL2_Mx9_1_Mx4_1_line3);
and3 M7_CSL2_Mx9_1_Mx4_1_Mux4_4(SumYbus_5, in4091, M7_CSL2_Mx9_1_Mx4_1_Not_ContLo, M7_CSL2_Mx9_1_Mx4_1_line4);
and3 M7_CSL2_Mx9_1_Mx4_1_Mux4_5(gnd, in4091, in4092, M7_CSL2_Mx9_1_Mx4_1_line5);
or4 M7_CSL2_Mx9_1_Mx4_1_Mux4_6(M7_CSL2_Mx9_1_Mx4_1_line2, M7_CSL2_Mx9_1_Mx4_1_line3, M7_CSL2_Mx9_1_Mx4_1_line4, M7_CSL2_Mx9_1_Mx4_1_line5, FYbus_5);
inv M7_CSL2_Mx9_1_Mx4_2_Mux4_0(in4092, M7_CSL2_Mx9_1_Mx4_2_Not_ContLo);
inv M7_CSL2_Mx9_1_Mx4_2_Mux4_1(in4091, M7_CSL2_Mx9_1_Mx4_2_Not_ContHi);
and3 M7_CSL2_Mx9_1_Mx4_2_Mux4_2(LogicYbus_6, M7_CSL2_Mx9_1_Mx4_2_Not_ContHi, M7_CSL2_Mx9_1_Mx4_2_Not_ContLo, M7_CSL2_Mx9_1_Mx4_2_line2);
and3 M7_CSL2_Mx9_1_Mx4_2_Mux4_3(in53, M7_CSL2_Mx9_1_Mx4_2_Not_ContHi, in4092, M7_CSL2_Mx9_1_Mx4_2_line3);
and3 M7_CSL2_Mx9_1_Mx4_2_Mux4_4(SumYbus_6, in4091, M7_CSL2_Mx9_1_Mx4_2_Not_ContLo, M7_CSL2_Mx9_1_Mx4_2_line4);
and3 M7_CSL2_Mx9_1_Mx4_2_Mux4_5(gnd, in4091, in4092, M7_CSL2_Mx9_1_Mx4_2_line5);
or4 M7_CSL2_Mx9_1_Mx4_2_Mux4_6(M7_CSL2_Mx9_1_Mx4_2_line2, M7_CSL2_Mx9_1_Mx4_2_line3, M7_CSL2_Mx9_1_Mx4_2_line4, M7_CSL2_Mx9_1_Mx4_2_line5, FYbus_6);
inv M7_CSL2_Mx9_1_Mx4_3_Mux4_0(in4092, M7_CSL2_Mx9_1_Mx4_3_Not_ContLo);
inv M7_CSL2_Mx9_1_Mx4_3_Mux4_1(in4091, M7_CSL2_Mx9_1_Mx4_3_Not_ContHi);
and3 M7_CSL2_Mx9_1_Mx4_3_Mux4_2(LogicYbus_7, M7_CSL2_Mx9_1_Mx4_3_Not_ContHi, M7_CSL2_Mx9_1_Mx4_3_Not_ContLo, M7_CSL2_Mx9_1_Mx4_3_line2);
and3 M7_CSL2_Mx9_1_Mx4_3_Mux4_3(in114, M7_CSL2_Mx9_1_Mx4_3_Not_ContHi, in4092, M7_CSL2_Mx9_1_Mx4_3_line3);
and3 M7_CSL2_Mx9_1_Mx4_3_Mux4_4(SumYbus_7, in4091, M7_CSL2_Mx9_1_Mx4_3_Not_ContLo, M7_CSL2_Mx9_1_Mx4_3_line4);
and3 M7_CSL2_Mx9_1_Mx4_3_Mux4_5(gnd, in4091, in4092, M7_CSL2_Mx9_1_Mx4_3_line5);
or4 M7_CSL2_Mx9_1_Mx4_3_Mux4_6(M7_CSL2_Mx9_1_Mx4_3_line2, M7_CSL2_Mx9_1_Mx4_3_line3, M7_CSL2_Mx9_1_Mx4_3_line4, M7_CSL2_Mx9_1_Mx4_3_line5, FYbus_7);
inv M7_CSL2_Mx9_2_Mux4_0(in4092, M7_CSL2_Mx9_2_Not_ContLo);
inv M7_CSL2_Mx9_2_Mux4_1(in4091, M7_CSL2_Mx9_2_Not_ContHi);
and3 M7_CSL2_Mx9_2_Mux4_2(LogicYbus_8, M7_CSL2_Mx9_2_Not_ContHi, M7_CSL2_Mx9_2_Not_ContLo, M7_CSL2_Mx9_2_line2);
and3 M7_CSL2_Mx9_2_Mux4_3(in115, M7_CSL2_Mx9_2_Not_ContHi, in4092, M7_CSL2_Mx9_2_line3);
and3 M7_CSL2_Mx9_2_Mux4_4(SumYbus_8, in4091, M7_CSL2_Mx9_2_Not_ContLo, M7_CSL2_Mx9_2_line4);
and3 M7_CSL2_Mx9_2_Mux4_5(gnd, in4091, in4092, M7_CSL2_Mx9_2_line5);
or4 M7_CSL2_Mx9_2_Mux4_6(M7_CSL2_Mx9_2_line2, M7_CSL2_Mx9_2_line3, M7_CSL2_Mx9_2_line4, M7_CSL2_Mx9_2_line5, FYbus_8);
inv M8_MF8_0_MF4_0_MXS0_Mux4_0(in1689, M8_MF8_0_MF4_0_MXS0_Not_ContLo);
inv M8_MF8_0_MF4_0_MXS0_Mux4_1(in1690, M8_MF8_0_MF4_0_MXS0_Not_ContHi);
and3 M8_MF8_0_MF4_0_MXS0_Mux4_2(FXbus_0, M8_MF8_0_MF4_0_MXS0_Not_ContHi, M8_MF8_0_MF4_0_MXS0_Not_ContLo, M8_MF8_0_MF4_0_MXS0_line2);
and3 M8_MF8_0_MF4_0_MXS0_Mux4_3(FYbus_0, M8_MF8_0_MF4_0_MXS0_Not_ContHi, in1689, M8_MF8_0_MF4_0_MXS0_line3);
and3 M8_MF8_0_MF4_0_MXS0_Mux4_4(in182, in1690, M8_MF8_0_MF4_0_MXS0_Not_ContLo, M8_MF8_0_MF4_0_MXS0_line4);
and3 M8_MF8_0_MF4_0_MXS0_Mux4_5(in185, in1690, in1689, M8_MF8_0_MF4_0_MXS0_line5);
or4 M8_MF8_0_MF4_0_MXS0_Mux4_6(M8_MF8_0_MF4_0_MXS0_line2, M8_MF8_0_MF4_0_MXS0_line3, M8_MF8_0_MF4_0_MXS0_line4, M8_MF8_0_MF4_0_MXS0_line5, M8_MF8_0_MF4_0_tempOut1);
inv M8_MF8_0_MF4_0_MXS1_Mux4_0(in1691, M8_MF8_0_MF4_0_MXS1_Not_ContLo);
inv M8_MF8_0_MF4_0_MXS1_Mux4_1(in1694, M8_MF8_0_MF4_0_MXS1_Not_ContHi);
and3 M8_MF8_0_MF4_0_MXS1_Mux4_2(FXbus_0, M8_MF8_0_MF4_0_MXS1_Not_ContHi, M8_MF8_0_MF4_0_MXS1_Not_ContLo, M8_MF8_0_MF4_0_MXS1_line2);
and3 M8_MF8_0_MF4_0_MXS1_Mux4_3(FYbus_0, M8_MF8_0_MF4_0_MXS1_Not_ContHi, in1691, M8_MF8_0_MF4_0_MXS1_line3);
and3 M8_MF8_0_MF4_0_MXS1_Mux4_4(in182, in1694, M8_MF8_0_MF4_0_MXS1_Not_ContLo, M8_MF8_0_MF4_0_MXS1_line4);
and3 M8_MF8_0_MF4_0_MXS1_Mux4_5(in185, in1694, in1691, M8_MF8_0_MF4_0_MXS1_line5);
or4 M8_MF8_0_MF4_0_MXS1_Mux4_6(M8_MF8_0_MF4_0_MXS1_line2, M8_MF8_0_MF4_0_MXS1_line3, M8_MF8_0_MF4_0_MXS1_line4, M8_MF8_0_MF4_0_MXS1_line5, M8_MF8_0_MF4_0_tempOut2);
inv M8_MF8_0_MF4_0_MXS2_Mux4_0(in4088, M8_MF8_0_MF4_0_MXS2_Not_ContLo);
inv M8_MF8_0_MF4_0_MXS2_Mux4_1(in4087, M8_MF8_0_MF4_0_MXS2_Not_ContHi);
and3 M8_MF8_0_MF4_0_MXS2_Mux4_2(FXbus_0, M8_MF8_0_MF4_0_MXS2_Not_ContHi, M8_MF8_0_MF4_0_MXS2_Not_ContLo, M8_MF8_0_MF4_0_MXS2_line2);
and3 M8_MF8_0_MF4_0_MXS2_Mux4_3(FYbus_0, M8_MF8_0_MF4_0_MXS2_Not_ContHi, in4088, M8_MF8_0_MF4_0_MXS2_line3);
and3 M8_MF8_0_MF4_0_MXS2_Mux4_4(in11, in4087, M8_MF8_0_MF4_0_MXS2_Not_ContLo, M8_MF8_0_MF4_0_MXS2_line4);
and3 M8_MF8_0_MF4_0_MXS2_Mux4_5(in61, in4087, in4088, M8_MF8_0_MF4_0_MXS2_line5);
or4 M8_MF8_0_MF4_0_MXS2_Mux4_6(M8_MF8_0_MF4_0_MXS2_line2, M8_MF8_0_MF4_0_MXS2_line3, M8_MF8_0_MF4_0_MXS2_line4, M8_MF8_0_MF4_0_MXS2_line5, out722);
inv M8_MF8_0_MF4_0_MXS3_Mux4_0(in4089, M8_MF8_0_MF4_0_MXS3_Not_ContLo);
inv M8_MF8_0_MF4_0_MXS3_Mux4_1(in4090, M8_MF8_0_MF4_0_MXS3_Not_ContHi);
and3 M8_MF8_0_MF4_0_MXS3_Mux4_2(FXbus_0, M8_MF8_0_MF4_0_MXS3_Not_ContHi, M8_MF8_0_MF4_0_MXS3_Not_ContLo, M8_MF8_0_MF4_0_MXS3_line2);
and3 M8_MF8_0_MF4_0_MXS3_Mux4_3(FYbus_0, M8_MF8_0_MF4_0_MXS3_Not_ContHi, in4089, M8_MF8_0_MF4_0_MXS3_line3);
and3 M8_MF8_0_MF4_0_MXS3_Mux4_4(in11, in4090, M8_MF8_0_MF4_0_MXS3_Not_ContLo, M8_MF8_0_MF4_0_MXS3_line4);
and3 M8_MF8_0_MF4_0_MXS3_Mux4_5(in61, in4090, in4089, M8_MF8_0_MF4_0_MXS3_line5);
or4 M8_MF8_0_MF4_0_MXS3_Mux4_6(M8_MF8_0_MF4_0_MXS3_line2, M8_MF8_0_MF4_0_MXS3_line3, M8_MF8_0_MF4_0_MXS3_line4, M8_MF8_0_MF4_0_MXS3_line5, out859);
and2 M8_MF8_0_MF4_0_MXS4(M8_MF8_0_MF4_0_tempOut1, in137, out661);
and2 M8_MF8_0_MF4_0_MXS5(M8_MF8_0_MF4_0_tempOut2, in137, out693);
inv M8_MF8_0_MF4_1_MXS0_Mux4_0(in1689, M8_MF8_0_MF4_1_MXS0_Not_ContLo);
inv M8_MF8_0_MF4_1_MXS0_Mux4_1(in1690, M8_MF8_0_MF4_1_MXS0_Not_ContHi);
and3 M8_MF8_0_MF4_1_MXS0_Mux4_2(FXbus_1, M8_MF8_0_MF4_1_MXS0_Not_ContHi, M8_MF8_0_MF4_1_MXS0_Not_ContLo, M8_MF8_0_MF4_1_MXS0_line2);
and3 M8_MF8_0_MF4_1_MXS0_Mux4_3(FYbus_1, M8_MF8_0_MF4_1_MXS0_Not_ContHi, in1689, M8_MF8_0_MF4_1_MXS0_line3);
and3 M8_MF8_0_MF4_1_MXS0_Mux4_4(in188, in1690, M8_MF8_0_MF4_1_MXS0_Not_ContLo, M8_MF8_0_MF4_1_MXS0_line4);
and3 M8_MF8_0_MF4_1_MXS0_Mux4_5(in158, in1690, in1689, M8_MF8_0_MF4_1_MXS0_line5);
or4 M8_MF8_0_MF4_1_MXS0_Mux4_6(M8_MF8_0_MF4_1_MXS0_line2, M8_MF8_0_MF4_1_MXS0_line3, M8_MF8_0_MF4_1_MXS0_line4, M8_MF8_0_MF4_1_MXS0_line5, M8_MF8_0_MF4_1_tempOut1);
inv M8_MF8_0_MF4_1_MXS1_Mux4_0(in1691, M8_MF8_0_MF4_1_MXS1_Not_ContLo);
inv M8_MF8_0_MF4_1_MXS1_Mux4_1(in1694, M8_MF8_0_MF4_1_MXS1_Not_ContHi);
and3 M8_MF8_0_MF4_1_MXS1_Mux4_2(FXbus_1, M8_MF8_0_MF4_1_MXS1_Not_ContHi, M8_MF8_0_MF4_1_MXS1_Not_ContLo, M8_MF8_0_MF4_1_MXS1_line2);
and3 M8_MF8_0_MF4_1_MXS1_Mux4_3(FYbus_1, M8_MF8_0_MF4_1_MXS1_Not_ContHi, in1691, M8_MF8_0_MF4_1_MXS1_line3);
and3 M8_MF8_0_MF4_1_MXS1_Mux4_4(in188, in1694, M8_MF8_0_MF4_1_MXS1_Not_ContLo, M8_MF8_0_MF4_1_MXS1_line4);
and3 M8_MF8_0_MF4_1_MXS1_Mux4_5(in158, in1694, in1691, M8_MF8_0_MF4_1_MXS1_line5);
or4 M8_MF8_0_MF4_1_MXS1_Mux4_6(M8_MF8_0_MF4_1_MXS1_line2, M8_MF8_0_MF4_1_MXS1_line3, M8_MF8_0_MF4_1_MXS1_line4, M8_MF8_0_MF4_1_MXS1_line5, M8_MF8_0_MF4_1_tempOut2);
inv M8_MF8_0_MF4_1_MXS2_Mux4_0(in4088, M8_MF8_0_MF4_1_MXS2_Not_ContLo);
inv M8_MF8_0_MF4_1_MXS2_Mux4_1(in4087, M8_MF8_0_MF4_1_MXS2_Not_ContHi);
and3 M8_MF8_0_MF4_1_MXS2_Mux4_2(FXbus_1, M8_MF8_0_MF4_1_MXS2_Not_ContHi, M8_MF8_0_MF4_1_MXS2_Not_ContLo, M8_MF8_0_MF4_1_MXS2_line2);
and3 M8_MF8_0_MF4_1_MXS2_Mux4_3(FYbus_1, M8_MF8_0_MF4_1_MXS2_Not_ContHi, in4088, M8_MF8_0_MF4_1_MXS2_line3);
and3 M8_MF8_0_MF4_1_MXS2_Mux4_4(in67, in4087, M8_MF8_0_MF4_1_MXS2_Not_ContLo, M8_MF8_0_MF4_1_MXS2_line4);
and3 M8_MF8_0_MF4_1_MXS2_Mux4_5(in70, in4087, in4088, M8_MF8_0_MF4_1_MXS2_line5);
or4 M8_MF8_0_MF4_1_MXS2_Mux4_6(M8_MF8_0_MF4_1_MXS2_line2, M8_MF8_0_MF4_1_MXS2_line3, M8_MF8_0_MF4_1_MXS2_line4, M8_MF8_0_MF4_1_MXS2_line5, out762);
inv M8_MF8_0_MF4_1_MXS3_Mux4_0(in4089, M8_MF8_0_MF4_1_MXS3_Not_ContLo);
inv M8_MF8_0_MF4_1_MXS3_Mux4_1(in4090, M8_MF8_0_MF4_1_MXS3_Not_ContHi);
and3 M8_MF8_0_MF4_1_MXS3_Mux4_2(FXbus_1, M8_MF8_0_MF4_1_MXS3_Not_ContHi, M8_MF8_0_MF4_1_MXS3_Not_ContLo, M8_MF8_0_MF4_1_MXS3_line2);
and3 M8_MF8_0_MF4_1_MXS3_Mux4_3(FYbus_1, M8_MF8_0_MF4_1_MXS3_Not_ContHi, in4089, M8_MF8_0_MF4_1_MXS3_line3);
and3 M8_MF8_0_MF4_1_MXS3_Mux4_4(in67, in4090, M8_MF8_0_MF4_1_MXS3_Not_ContLo, M8_MF8_0_MF4_1_MXS3_line4);
and3 M8_MF8_0_MF4_1_MXS3_Mux4_5(in70, in4090, in4089, M8_MF8_0_MF4_1_MXS3_line5);
or4 M8_MF8_0_MF4_1_MXS3_Mux4_6(M8_MF8_0_MF4_1_MXS3_line2, M8_MF8_0_MF4_1_MXS3_line3, M8_MF8_0_MF4_1_MXS3_line4, M8_MF8_0_MF4_1_MXS3_line5, out802);
and2 M8_MF8_0_MF4_1_MXS4(M8_MF8_0_MF4_1_tempOut1, in137, out664);
and2 M8_MF8_0_MF4_1_MXS5(M8_MF8_0_MF4_1_tempOut2, in137, out696);
inv M8_MF8_0_MF4_2_MXS0_Mux4_0(in1689, M8_MF8_0_MF4_2_MXS0_Not_ContLo);
inv M8_MF8_0_MF4_2_MXS0_Mux4_1(in1690, M8_MF8_0_MF4_2_MXS0_Not_ContHi);
and3 M8_MF8_0_MF4_2_MXS0_Mux4_2(FXbus_2, M8_MF8_0_MF4_2_MXS0_Not_ContHi, M8_MF8_0_MF4_2_MXS0_Not_ContLo, M8_MF8_0_MF4_2_MXS0_line2);
and3 M8_MF8_0_MF4_2_MXS0_Mux4_3(FYbus_2, M8_MF8_0_MF4_2_MXS0_Not_ContHi, in1689, M8_MF8_0_MF4_2_MXS0_line3);
and3 M8_MF8_0_MF4_2_MXS0_Mux4_4(in155, in1690, M8_MF8_0_MF4_2_MXS0_Not_ContLo, M8_MF8_0_MF4_2_MXS0_line4);
and3 M8_MF8_0_MF4_2_MXS0_Mux4_5(in152, in1690, in1689, M8_MF8_0_MF4_2_MXS0_line5);
or4 M8_MF8_0_MF4_2_MXS0_Mux4_6(M8_MF8_0_MF4_2_MXS0_line2, M8_MF8_0_MF4_2_MXS0_line3, M8_MF8_0_MF4_2_MXS0_line4, M8_MF8_0_MF4_2_MXS0_line5, M8_MF8_0_MF4_2_tempOut1);
inv M8_MF8_0_MF4_2_MXS1_Mux4_0(in1691, M8_MF8_0_MF4_2_MXS1_Not_ContLo);
inv M8_MF8_0_MF4_2_MXS1_Mux4_1(in1694, M8_MF8_0_MF4_2_MXS1_Not_ContHi);
and3 M8_MF8_0_MF4_2_MXS1_Mux4_2(FXbus_2, M8_MF8_0_MF4_2_MXS1_Not_ContHi, M8_MF8_0_MF4_2_MXS1_Not_ContLo, M8_MF8_0_MF4_2_MXS1_line2);
and3 M8_MF8_0_MF4_2_MXS1_Mux4_3(FYbus_2, M8_MF8_0_MF4_2_MXS1_Not_ContHi, in1691, M8_MF8_0_MF4_2_MXS1_line3);
and3 M8_MF8_0_MF4_2_MXS1_Mux4_4(in155, in1694, M8_MF8_0_MF4_2_MXS1_Not_ContLo, M8_MF8_0_MF4_2_MXS1_line4);
and3 M8_MF8_0_MF4_2_MXS1_Mux4_5(in152, in1694, in1691, M8_MF8_0_MF4_2_MXS1_line5);
or4 M8_MF8_0_MF4_2_MXS1_Mux4_6(M8_MF8_0_MF4_2_MXS1_line2, M8_MF8_0_MF4_2_MXS1_line3, M8_MF8_0_MF4_2_MXS1_line4, M8_MF8_0_MF4_2_MXS1_line5, M8_MF8_0_MF4_2_tempOut2);
inv M8_MF8_0_MF4_2_MXS2_Mux4_0(in4088, M8_MF8_0_MF4_2_MXS2_Not_ContLo);
inv M8_MF8_0_MF4_2_MXS2_Mux4_1(in4087, M8_MF8_0_MF4_2_MXS2_Not_ContHi);
and3 M8_MF8_0_MF4_2_MXS2_Mux4_2(FXbus_2, M8_MF8_0_MF4_2_MXS2_Not_ContHi, M8_MF8_0_MF4_2_MXS2_Not_ContLo, M8_MF8_0_MF4_2_MXS2_line2);
and3 M8_MF8_0_MF4_2_MXS2_Mux4_3(FYbus_2, M8_MF8_0_MF4_2_MXS2_Not_ContHi, in4088, M8_MF8_0_MF4_2_MXS2_line3);
and3 M8_MF8_0_MF4_2_MXS2_Mux4_4(in73, in4087, M8_MF8_0_MF4_2_MXS2_Not_ContLo, M8_MF8_0_MF4_2_MXS2_line4);
and3 M8_MF8_0_MF4_2_MXS2_Mux4_5(in17, in4087, in4088, M8_MF8_0_MF4_2_MXS2_line5);
or4 M8_MF8_0_MF4_2_MXS2_Mux4_6(M8_MF8_0_MF4_2_MXS2_line2, M8_MF8_0_MF4_2_MXS2_line3, M8_MF8_0_MF4_2_MXS2_line4, M8_MF8_0_MF4_2_MXS2_line5, out757);
inv M8_MF8_0_MF4_2_MXS3_Mux4_0(in4089, M8_MF8_0_MF4_2_MXS3_Not_ContLo);
inv M8_MF8_0_MF4_2_MXS3_Mux4_1(in4090, M8_MF8_0_MF4_2_MXS3_Not_ContHi);
and3 M8_MF8_0_MF4_2_MXS3_Mux4_2(FXbus_2, M8_MF8_0_MF4_2_MXS3_Not_ContHi, M8_MF8_0_MF4_2_MXS3_Not_ContLo, M8_MF8_0_MF4_2_MXS3_line2);
and3 M8_MF8_0_MF4_2_MXS3_Mux4_3(FYbus_2, M8_MF8_0_MF4_2_MXS3_Not_ContHi, in4089, M8_MF8_0_MF4_2_MXS3_line3);
and3 M8_MF8_0_MF4_2_MXS3_Mux4_4(in73, in4090, M8_MF8_0_MF4_2_MXS3_Not_ContLo, M8_MF8_0_MF4_2_MXS3_line4);
and3 M8_MF8_0_MF4_2_MXS3_Mux4_5(in17, in4090, in4089, M8_MF8_0_MF4_2_MXS3_line5);
or4 M8_MF8_0_MF4_2_MXS3_Mux4_6(M8_MF8_0_MF4_2_MXS3_line2, M8_MF8_0_MF4_2_MXS3_line3, M8_MF8_0_MF4_2_MXS3_line4, M8_MF8_0_MF4_2_MXS3_line5, out797);
and2 M8_MF8_0_MF4_2_MXS4(M8_MF8_0_MF4_2_tempOut1, in137, out667);
and2 M8_MF8_0_MF4_2_MXS5(M8_MF8_0_MF4_2_tempOut2, in137, out699);
inv M8_MF8_0_MF8_3_MXS0_Mux4_0(in1689, M8_MF8_0_MF8_3_MXS0_Not_ContLo);
inv M8_MF8_0_MF8_3_MXS0_Mux4_1(in1690, M8_MF8_0_MF8_3_MXS0_Not_ContHi);
and3 M8_MF8_0_MF8_3_MXS0_Mux4_2(FXbus_3, M8_MF8_0_MF8_3_MXS0_Not_ContHi, M8_MF8_0_MF8_3_MXS0_Not_ContLo, M8_MF8_0_MF8_3_MXS0_line2);
and3 M8_MF8_0_MF8_3_MXS0_Mux4_3(FYbus_3, M8_MF8_0_MF8_3_MXS0_Not_ContHi, in1689, M8_MF8_0_MF8_3_MXS0_line3);
and3 M8_MF8_0_MF8_3_MXS0_Mux4_4(in149, in1690, M8_MF8_0_MF8_3_MXS0_Not_ContLo, M8_MF8_0_MF8_3_MXS0_line4);
and3 M8_MF8_0_MF8_3_MXS0_Mux4_5(in146, in1690, in1689, M8_MF8_0_MF8_3_MXS0_line5);
or4 M8_MF8_0_MF8_3_MXS0_Mux4_6(M8_MF8_0_MF8_3_MXS0_line2, M8_MF8_0_MF8_3_MXS0_line3, M8_MF8_0_MF8_3_MXS0_line4, M8_MF8_0_MF8_3_MXS0_line5, M8_MF8_0_MF8_3_tempOut1);
inv M8_MF8_0_MF8_3_MXS1_Mux4_0(in1691, M8_MF8_0_MF8_3_MXS1_Not_ContLo);
inv M8_MF8_0_MF8_3_MXS1_Mux4_1(in1694, M8_MF8_0_MF8_3_MXS1_Not_ContHi);
and3 M8_MF8_0_MF8_3_MXS1_Mux4_2(FXbus_3, M8_MF8_0_MF8_3_MXS1_Not_ContHi, M8_MF8_0_MF8_3_MXS1_Not_ContLo, M8_MF8_0_MF8_3_MXS1_line2);
and3 M8_MF8_0_MF8_3_MXS1_Mux4_3(FYbus_3, M8_MF8_0_MF8_3_MXS1_Not_ContHi, in1691, M8_MF8_0_MF8_3_MXS1_line3);
and3 M8_MF8_0_MF8_3_MXS1_Mux4_4(in149, in1694, M8_MF8_0_MF8_3_MXS1_Not_ContLo, M8_MF8_0_MF8_3_MXS1_line4);
and3 M8_MF8_0_MF8_3_MXS1_Mux4_5(in146, in1694, in1691, M8_MF8_0_MF8_3_MXS1_line5);
or4 M8_MF8_0_MF8_3_MXS1_Mux4_6(M8_MF8_0_MF8_3_MXS1_line2, M8_MF8_0_MF8_3_MXS1_line3, M8_MF8_0_MF8_3_MXS1_line4, M8_MF8_0_MF8_3_MXS1_line5, M8_MF8_0_MF8_3_tempOut2);
inv M8_MF8_0_MF8_3_MXS2_Mux4_0(in4088, M8_MF8_0_MF8_3_MXS2_Not_ContLo);
inv M8_MF8_0_MF8_3_MXS2_Mux4_1(in4087, M8_MF8_0_MF8_3_MXS2_Not_ContHi);
and3 M8_MF8_0_MF8_3_MXS2_Mux4_2(FXbus_3, M8_MF8_0_MF8_3_MXS2_Not_ContHi, M8_MF8_0_MF8_3_MXS2_Not_ContLo, M8_MF8_0_MF8_3_MXS2_line2);
and3 M8_MF8_0_MF8_3_MXS2_Mux4_3(FYbus_3, M8_MF8_0_MF8_3_MXS2_Not_ContHi, in4088, M8_MF8_0_MF8_3_MXS2_line3);
and3 M8_MF8_0_MF8_3_MXS2_Mux4_4(in76, in4087, M8_MF8_0_MF8_3_MXS2_Not_ContLo, M8_MF8_0_MF8_3_MXS2_line4);
and3 M8_MF8_0_MF8_3_MXS2_Mux4_5(in20, in4087, in4088, M8_MF8_0_MF8_3_MXS2_line5);
or4 M8_MF8_0_MF8_3_MXS2_Mux4_6(M8_MF8_0_MF8_3_MXS2_line2, M8_MF8_0_MF8_3_MXS2_line3, M8_MF8_0_MF8_3_MXS2_line4, M8_MF8_0_MF8_3_MXS2_line5, out752);
inv M8_MF8_0_MF8_3_MXS3_Mux4_0(in4089, M8_MF8_0_MF8_3_MXS3_Not_ContLo);
inv M8_MF8_0_MF8_3_MXS3_Mux4_1(in4090, M8_MF8_0_MF8_3_MXS3_Not_ContHi);
and3 M8_MF8_0_MF8_3_MXS3_Mux4_2(FXbus_3, M8_MF8_0_MF8_3_MXS3_Not_ContHi, M8_MF8_0_MF8_3_MXS3_Not_ContLo, M8_MF8_0_MF8_3_MXS3_line2);
and3 M8_MF8_0_MF8_3_MXS3_Mux4_3(FYbus_3, M8_MF8_0_MF8_3_MXS3_Not_ContHi, in4089, M8_MF8_0_MF8_3_MXS3_line3);
and3 M8_MF8_0_MF8_3_MXS3_Mux4_4(in76, in4090, M8_MF8_0_MF8_3_MXS3_Not_ContLo, M8_MF8_0_MF8_3_MXS3_line4);
and3 M8_MF8_0_MF8_3_MXS3_Mux4_5(in20, in4090, in4089, M8_MF8_0_MF8_3_MXS3_line5);
or4 M8_MF8_0_MF8_3_MXS3_Mux4_6(M8_MF8_0_MF8_3_MXS3_line2, M8_MF8_0_MF8_3_MXS3_line3, M8_MF8_0_MF8_3_MXS3_line4, M8_MF8_0_MF8_3_MXS3_line5, out792);
and2 M8_MF8_0_MF8_3_MXS4(M8_MF8_0_MF8_3_tempOut1, in137, out670);
and2 M8_MF8_0_MF8_3_MXS5(M8_MF8_0_MF8_3_tempOut2, in137, out702);
inv M8_MF8_1_MF4_0_MXS0_Mux4_0(in1689, M8_MF8_1_MF4_0_MXS0_Not_ContLo);
inv M8_MF8_1_MF4_0_MXS0_Mux4_1(in1690, M8_MF8_1_MF4_0_MXS0_Not_ContHi);
and3 M8_MF8_1_MF4_0_MXS0_Mux4_2(FXbus_4, M8_MF8_1_MF4_0_MXS0_Not_ContHi, M8_MF8_1_MF4_0_MXS0_Not_ContLo, M8_MF8_1_MF4_0_MXS0_line2);
and3 M8_MF8_1_MF4_0_MXS0_Mux4_3(FYbus_4, M8_MF8_1_MF4_0_MXS0_Not_ContHi, in1689, M8_MF8_1_MF4_0_MXS0_line3);
and3 M8_MF8_1_MF4_0_MXS0_Mux4_4(in200, in1690, M8_MF8_1_MF4_0_MXS0_Not_ContLo, M8_MF8_1_MF4_0_MXS0_line4);
and3 M8_MF8_1_MF4_0_MXS0_Mux4_5(in170, in1690, in1689, M8_MF8_1_MF4_0_MXS0_line5);
or4 M8_MF8_1_MF4_0_MXS0_Mux4_6(M8_MF8_1_MF4_0_MXS0_line2, M8_MF8_1_MF4_0_MXS0_line3, M8_MF8_1_MF4_0_MXS0_line4, M8_MF8_1_MF4_0_MXS0_line5, M8_MF8_1_MF4_0_tempOut1);
inv M8_MF8_1_MF4_0_MXS1_Mux4_0(in1691, M8_MF8_1_MF4_0_MXS1_Not_ContLo);
inv M8_MF8_1_MF4_0_MXS1_Mux4_1(in1694, M8_MF8_1_MF4_0_MXS1_Not_ContHi);
and3 M8_MF8_1_MF4_0_MXS1_Mux4_2(FXbus_4, M8_MF8_1_MF4_0_MXS1_Not_ContHi, M8_MF8_1_MF4_0_MXS1_Not_ContLo, M8_MF8_1_MF4_0_MXS1_line2);
and3 M8_MF8_1_MF4_0_MXS1_Mux4_3(FYbus_4, M8_MF8_1_MF4_0_MXS1_Not_ContHi, in1691, M8_MF8_1_MF4_0_MXS1_line3);
and3 M8_MF8_1_MF4_0_MXS1_Mux4_4(in200, in1694, M8_MF8_1_MF4_0_MXS1_Not_ContLo, M8_MF8_1_MF4_0_MXS1_line4);
and3 M8_MF8_1_MF4_0_MXS1_Mux4_5(in170, in1694, in1691, M8_MF8_1_MF4_0_MXS1_line5);
or4 M8_MF8_1_MF4_0_MXS1_Mux4_6(M8_MF8_1_MF4_0_MXS1_line2, M8_MF8_1_MF4_0_MXS1_line3, M8_MF8_1_MF4_0_MXS1_line4, M8_MF8_1_MF4_0_MXS1_line5, M8_MF8_1_MF4_0_tempOut2);
inv M8_MF8_1_MF4_0_MXS2_Mux4_0(in4088, M8_MF8_1_MF4_0_MXS2_Not_ContLo);
inv M8_MF8_1_MF4_0_MXS2_Mux4_1(in4087, M8_MF8_1_MF4_0_MXS2_Not_ContHi);
and3 M8_MF8_1_MF4_0_MXS2_Mux4_2(FXbus_4, M8_MF8_1_MF4_0_MXS2_Not_ContHi, M8_MF8_1_MF4_0_MXS2_Not_ContLo, M8_MF8_1_MF4_0_MXS2_line2);
and3 M8_MF8_1_MF4_0_MXS2_Mux4_3(FYbus_4, M8_MF8_1_MF4_0_MXS2_Not_ContHi, in4088, M8_MF8_1_MF4_0_MXS2_line3);
and3 M8_MF8_1_MF4_0_MXS2_Mux4_4(in43, in4087, M8_MF8_1_MF4_0_MXS2_Not_ContLo, M8_MF8_1_MF4_0_MXS2_line4);
and3 M8_MF8_1_MF4_0_MXS2_Mux4_5(in37, in4087, in4088, M8_MF8_1_MF4_0_MXS2_line5);
or4 M8_MF8_1_MF4_0_MXS2_Mux4_6(M8_MF8_1_MF4_0_MXS2_line2, M8_MF8_1_MF4_0_MXS2_line3, M8_MF8_1_MF4_0_MXS2_line4, M8_MF8_1_MF4_0_MXS2_line5, out747);
inv M8_MF8_1_MF4_0_MXS3_Mux4_0(in4089, M8_MF8_1_MF4_0_MXS3_Not_ContLo);
inv M8_MF8_1_MF4_0_MXS3_Mux4_1(in4090, M8_MF8_1_MF4_0_MXS3_Not_ContHi);
and3 M8_MF8_1_MF4_0_MXS3_Mux4_2(FXbus_4, M8_MF8_1_MF4_0_MXS3_Not_ContHi, M8_MF8_1_MF4_0_MXS3_Not_ContLo, M8_MF8_1_MF4_0_MXS3_line2);
and3 M8_MF8_1_MF4_0_MXS3_Mux4_3(FYbus_4, M8_MF8_1_MF4_0_MXS3_Not_ContHi, in4089, M8_MF8_1_MF4_0_MXS3_line3);
and3 M8_MF8_1_MF4_0_MXS3_Mux4_4(in43, in4090, M8_MF8_1_MF4_0_MXS3_Not_ContLo, M8_MF8_1_MF4_0_MXS3_line4);
and3 M8_MF8_1_MF4_0_MXS3_Mux4_5(in37, in4090, in4089, M8_MF8_1_MF4_0_MXS3_line5);
or4 M8_MF8_1_MF4_0_MXS3_Mux4_6(M8_MF8_1_MF4_0_MXS3_line2, M8_MF8_1_MF4_0_MXS3_line3, M8_MF8_1_MF4_0_MXS3_line4, M8_MF8_1_MF4_0_MXS3_line5, out787);
and2 M8_MF8_1_MF4_0_MXS4(M8_MF8_1_MF4_0_tempOut1, in137, out642);
and2 M8_MF8_1_MF4_0_MXS5(M8_MF8_1_MF4_0_tempOut2, in137, out676);
inv M8_MF8_1_MF4_1_MXS0_Mux4_0(in1689, M8_MF8_1_MF4_1_MXS0_Not_ContLo);
inv M8_MF8_1_MF4_1_MXS0_Mux4_1(in1690, M8_MF8_1_MF4_1_MXS0_Not_ContHi);
and3 M8_MF8_1_MF4_1_MXS0_Mux4_2(FXbus_5, M8_MF8_1_MF4_1_MXS0_Not_ContHi, M8_MF8_1_MF4_1_MXS0_Not_ContLo, M8_MF8_1_MF4_1_MXS0_line2);
and3 M8_MF8_1_MF4_1_MXS0_Mux4_3(FYbus_5, M8_MF8_1_MF4_1_MXS0_Not_ContHi, in1689, M8_MF8_1_MF4_1_MXS0_line3);
and3 M8_MF8_1_MF4_1_MXS0_Mux4_4(in203, in1690, M8_MF8_1_MF4_1_MXS0_Not_ContLo, M8_MF8_1_MF4_1_MXS0_line4);
and3 M8_MF8_1_MF4_1_MXS0_Mux4_5(in173, in1690, in1689, M8_MF8_1_MF4_1_MXS0_line5);
or4 M8_MF8_1_MF4_1_MXS0_Mux4_6(M8_MF8_1_MF4_1_MXS0_line2, M8_MF8_1_MF4_1_MXS0_line3, M8_MF8_1_MF4_1_MXS0_line4, M8_MF8_1_MF4_1_MXS0_line5, M8_MF8_1_MF4_1_tempOut1);
inv M8_MF8_1_MF4_1_MXS1_Mux4_0(in1691, M8_MF8_1_MF4_1_MXS1_Not_ContLo);
inv M8_MF8_1_MF4_1_MXS1_Mux4_1(in1694, M8_MF8_1_MF4_1_MXS1_Not_ContHi);
and3 M8_MF8_1_MF4_1_MXS1_Mux4_2(FXbus_5, M8_MF8_1_MF4_1_MXS1_Not_ContHi, M8_MF8_1_MF4_1_MXS1_Not_ContLo, M8_MF8_1_MF4_1_MXS1_line2);
and3 M8_MF8_1_MF4_1_MXS1_Mux4_3(FYbus_5, M8_MF8_1_MF4_1_MXS1_Not_ContHi, in1691, M8_MF8_1_MF4_1_MXS1_line3);
and3 M8_MF8_1_MF4_1_MXS1_Mux4_4(in203, in1694, M8_MF8_1_MF4_1_MXS1_Not_ContLo, M8_MF8_1_MF4_1_MXS1_line4);
and3 M8_MF8_1_MF4_1_MXS1_Mux4_5(in173, in1694, in1691, M8_MF8_1_MF4_1_MXS1_line5);
or4 M8_MF8_1_MF4_1_MXS1_Mux4_6(M8_MF8_1_MF4_1_MXS1_line2, M8_MF8_1_MF4_1_MXS1_line3, M8_MF8_1_MF4_1_MXS1_line4, M8_MF8_1_MF4_1_MXS1_line5, M8_MF8_1_MF4_1_tempOut2);
inv M8_MF8_1_MF4_1_MXS2_Mux4_0(in4088, M8_MF8_1_MF4_1_MXS2_Not_ContLo);
inv M8_MF8_1_MF4_1_MXS2_Mux4_1(in4087, M8_MF8_1_MF4_1_MXS2_Not_ContHi);
and3 M8_MF8_1_MF4_1_MXS2_Mux4_2(FXbus_5, M8_MF8_1_MF4_1_MXS2_Not_ContHi, M8_MF8_1_MF4_1_MXS2_Not_ContLo, M8_MF8_1_MF4_1_MXS2_line2);
and3 M8_MF8_1_MF4_1_MXS2_Mux4_3(FYbus_5, M8_MF8_1_MF4_1_MXS2_Not_ContHi, in4088, M8_MF8_1_MF4_1_MXS2_line3);
and3 M8_MF8_1_MF4_1_MXS2_Mux4_4(in91, in4087, M8_MF8_1_MF4_1_MXS2_Not_ContLo, M8_MF8_1_MF4_1_MXS2_line4);
and3 M8_MF8_1_MF4_1_MXS2_Mux4_5(in40, in4087, in4088, M8_MF8_1_MF4_1_MXS2_line5);
or4 M8_MF8_1_MF4_1_MXS2_Mux4_6(M8_MF8_1_MF4_1_MXS2_line2, M8_MF8_1_MF4_1_MXS2_line3, M8_MF8_1_MF4_1_MXS2_line4, M8_MF8_1_MF4_1_MXS2_line5, out742);
inv M8_MF8_1_MF4_1_MXS3_Mux4_0(in4089, M8_MF8_1_MF4_1_MXS3_Not_ContLo);
inv M8_MF8_1_MF4_1_MXS3_Mux4_1(in4090, M8_MF8_1_MF4_1_MXS3_Not_ContHi);
and3 M8_MF8_1_MF4_1_MXS3_Mux4_2(FXbus_5, M8_MF8_1_MF4_1_MXS3_Not_ContHi, M8_MF8_1_MF4_1_MXS3_Not_ContLo, M8_MF8_1_MF4_1_MXS3_line2);
and3 M8_MF8_1_MF4_1_MXS3_Mux4_3(FYbus_5, M8_MF8_1_MF4_1_MXS3_Not_ContHi, in4089, M8_MF8_1_MF4_1_MXS3_line3);
and3 M8_MF8_1_MF4_1_MXS3_Mux4_4(in91, in4090, M8_MF8_1_MF4_1_MXS3_Not_ContLo, M8_MF8_1_MF4_1_MXS3_line4);
and3 M8_MF8_1_MF4_1_MXS3_Mux4_5(in40, in4090, in4089, M8_MF8_1_MF4_1_MXS3_line5);
or4 M8_MF8_1_MF4_1_MXS3_Mux4_6(M8_MF8_1_MF4_1_MXS3_line2, M8_MF8_1_MF4_1_MXS3_line3, M8_MF8_1_MF4_1_MXS3_line4, M8_MF8_1_MF4_1_MXS3_line5, out782);
and2 M8_MF8_1_MF4_1_MXS4(M8_MF8_1_MF4_1_tempOut1, in137, out645);
and2 M8_MF8_1_MF4_1_MXS5(M8_MF8_1_MF4_1_tempOut2, in137, out679);
inv M8_MF8_1_MF4_2_MXS0_Mux4_0(in1689, M8_MF8_1_MF4_2_MXS0_Not_ContLo);
inv M8_MF8_1_MF4_2_MXS0_Mux4_1(in1690, M8_MF8_1_MF4_2_MXS0_Not_ContHi);
and3 M8_MF8_1_MF4_2_MXS0_Mux4_2(FXbus_6, M8_MF8_1_MF4_2_MXS0_Not_ContHi, M8_MF8_1_MF4_2_MXS0_Not_ContLo, M8_MF8_1_MF4_2_MXS0_line2);
and3 M8_MF8_1_MF4_2_MXS0_Mux4_3(FYbus_6, M8_MF8_1_MF4_2_MXS0_Not_ContHi, in1689, M8_MF8_1_MF4_2_MXS0_line3);
and3 M8_MF8_1_MF4_2_MXS0_Mux4_4(in197, in1690, M8_MF8_1_MF4_2_MXS0_Not_ContLo, M8_MF8_1_MF4_2_MXS0_line4);
and3 M8_MF8_1_MF4_2_MXS0_Mux4_5(in167, in1690, in1689, M8_MF8_1_MF4_2_MXS0_line5);
or4 M8_MF8_1_MF4_2_MXS0_Mux4_6(M8_MF8_1_MF4_2_MXS0_line2, M8_MF8_1_MF4_2_MXS0_line3, M8_MF8_1_MF4_2_MXS0_line4, M8_MF8_1_MF4_2_MXS0_line5, M8_MF8_1_MF4_2_tempOut1);
inv M8_MF8_1_MF4_2_MXS1_Mux4_0(in1691, M8_MF8_1_MF4_2_MXS1_Not_ContLo);
inv M8_MF8_1_MF4_2_MXS1_Mux4_1(in1694, M8_MF8_1_MF4_2_MXS1_Not_ContHi);
and3 M8_MF8_1_MF4_2_MXS1_Mux4_2(FXbus_6, M8_MF8_1_MF4_2_MXS1_Not_ContHi, M8_MF8_1_MF4_2_MXS1_Not_ContLo, M8_MF8_1_MF4_2_MXS1_line2);
and3 M8_MF8_1_MF4_2_MXS1_Mux4_3(FYbus_6, M8_MF8_1_MF4_2_MXS1_Not_ContHi, in1691, M8_MF8_1_MF4_2_MXS1_line3);
and3 M8_MF8_1_MF4_2_MXS1_Mux4_4(in197, in1694, M8_MF8_1_MF4_2_MXS1_Not_ContLo, M8_MF8_1_MF4_2_MXS1_line4);
and3 M8_MF8_1_MF4_2_MXS1_Mux4_5(in167, in1694, in1691, M8_MF8_1_MF4_2_MXS1_line5);
or4 M8_MF8_1_MF4_2_MXS1_Mux4_6(M8_MF8_1_MF4_2_MXS1_line2, M8_MF8_1_MF4_2_MXS1_line3, M8_MF8_1_MF4_2_MXS1_line4, M8_MF8_1_MF4_2_MXS1_line5, M8_MF8_1_MF4_2_tempOut2);
inv M8_MF8_1_MF4_2_MXS2_Mux4_0(in4088, M8_MF8_1_MF4_2_MXS2_Not_ContLo);
inv M8_MF8_1_MF4_2_MXS2_Mux4_1(in4087, M8_MF8_1_MF4_2_MXS2_Not_ContHi);
and3 M8_MF8_1_MF4_2_MXS2_Mux4_2(FXbus_6, M8_MF8_1_MF4_2_MXS2_Not_ContHi, M8_MF8_1_MF4_2_MXS2_Not_ContLo, M8_MF8_1_MF4_2_MXS2_line2);
and3 M8_MF8_1_MF4_2_MXS2_Mux4_3(FYbus_6, M8_MF8_1_MF4_2_MXS2_Not_ContHi, in4088, M8_MF8_1_MF4_2_MXS2_line3);
and3 M8_MF8_1_MF4_2_MXS2_Mux4_4(in100, in4087, M8_MF8_1_MF4_2_MXS2_Not_ContLo, M8_MF8_1_MF4_2_MXS2_line4);
and3 M8_MF8_1_MF4_2_MXS2_Mux4_5(in103, in4087, in4088, M8_MF8_1_MF4_2_MXS2_line5);
or4 M8_MF8_1_MF4_2_MXS2_Mux4_6(M8_MF8_1_MF4_2_MXS2_line2, M8_MF8_1_MF4_2_MXS2_line3, M8_MF8_1_MF4_2_MXS2_line4, M8_MF8_1_MF4_2_MXS2_line5, out737);
inv M8_MF8_1_MF4_2_MXS3_Mux4_0(in4089, M8_MF8_1_MF4_2_MXS3_Not_ContLo);
inv M8_MF8_1_MF4_2_MXS3_Mux4_1(in4090, M8_MF8_1_MF4_2_MXS3_Not_ContHi);
and3 M8_MF8_1_MF4_2_MXS3_Mux4_2(FXbus_6, M8_MF8_1_MF4_2_MXS3_Not_ContHi, M8_MF8_1_MF4_2_MXS3_Not_ContLo, M8_MF8_1_MF4_2_MXS3_line2);
and3 M8_MF8_1_MF4_2_MXS3_Mux4_3(FYbus_6, M8_MF8_1_MF4_2_MXS3_Not_ContHi, in4089, M8_MF8_1_MF4_2_MXS3_line3);
and3 M8_MF8_1_MF4_2_MXS3_Mux4_4(in100, in4090, M8_MF8_1_MF4_2_MXS3_Not_ContLo, M8_MF8_1_MF4_2_MXS3_line4);
and3 M8_MF8_1_MF4_2_MXS3_Mux4_5(in103, in4090, in4089, M8_MF8_1_MF4_2_MXS3_line5);
or4 M8_MF8_1_MF4_2_MXS3_Mux4_6(M8_MF8_1_MF4_2_MXS3_line2, M8_MF8_1_MF4_2_MXS3_line3, M8_MF8_1_MF4_2_MXS3_line4, M8_MF8_1_MF4_2_MXS3_line5, out777);
and2 M8_MF8_1_MF4_2_MXS4(M8_MF8_1_MF4_2_tempOut1, in137, out648);
and2 M8_MF8_1_MF4_2_MXS5(M8_MF8_1_MF4_2_tempOut2, in137, out682);
inv M8_MF8_1_MF8_3_MXS0_Mux4_0(in1689, M8_MF8_1_MF8_3_MXS0_Not_ContLo);
inv M8_MF8_1_MF8_3_MXS0_Mux4_1(in1690, M8_MF8_1_MF8_3_MXS0_Not_ContHi);
and3 M8_MF8_1_MF8_3_MXS0_Mux4_2(FXbus_7, M8_MF8_1_MF8_3_MXS0_Not_ContHi, M8_MF8_1_MF8_3_MXS0_Not_ContLo, M8_MF8_1_MF8_3_MXS0_line2);
and3 M8_MF8_1_MF8_3_MXS0_Mux4_3(FYbus_7, M8_MF8_1_MF8_3_MXS0_Not_ContHi, in1689, M8_MF8_1_MF8_3_MXS0_line3);
and3 M8_MF8_1_MF8_3_MXS0_Mux4_4(in194, in1690, M8_MF8_1_MF8_3_MXS0_Not_ContLo, M8_MF8_1_MF8_3_MXS0_line4);
and3 M8_MF8_1_MF8_3_MXS0_Mux4_5(in164, in1690, in1689, M8_MF8_1_MF8_3_MXS0_line5);
or4 M8_MF8_1_MF8_3_MXS0_Mux4_6(M8_MF8_1_MF8_3_MXS0_line2, M8_MF8_1_MF8_3_MXS0_line3, M8_MF8_1_MF8_3_MXS0_line4, M8_MF8_1_MF8_3_MXS0_line5, M8_MF8_1_MF8_3_tempOut1);
inv M8_MF8_1_MF8_3_MXS1_Mux4_0(in1691, M8_MF8_1_MF8_3_MXS1_Not_ContLo);
inv M8_MF8_1_MF8_3_MXS1_Mux4_1(in1694, M8_MF8_1_MF8_3_MXS1_Not_ContHi);
and3 M8_MF8_1_MF8_3_MXS1_Mux4_2(FXbus_7, M8_MF8_1_MF8_3_MXS1_Not_ContHi, M8_MF8_1_MF8_3_MXS1_Not_ContLo, M8_MF8_1_MF8_3_MXS1_line2);
and3 M8_MF8_1_MF8_3_MXS1_Mux4_3(FYbus_7, M8_MF8_1_MF8_3_MXS1_Not_ContHi, in1691, M8_MF8_1_MF8_3_MXS1_line3);
and3 M8_MF8_1_MF8_3_MXS1_Mux4_4(in194, in1694, M8_MF8_1_MF8_3_MXS1_Not_ContLo, M8_MF8_1_MF8_3_MXS1_line4);
and3 M8_MF8_1_MF8_3_MXS1_Mux4_5(in164, in1694, in1691, M8_MF8_1_MF8_3_MXS1_line5);
or4 M8_MF8_1_MF8_3_MXS1_Mux4_6(M8_MF8_1_MF8_3_MXS1_line2, M8_MF8_1_MF8_3_MXS1_line3, M8_MF8_1_MF8_3_MXS1_line4, M8_MF8_1_MF8_3_MXS1_line5, M8_MF8_1_MF8_3_tempOut2);
inv M8_MF8_1_MF8_3_MXS2_Mux4_0(in4088, M8_MF8_1_MF8_3_MXS2_Not_ContLo);
inv M8_MF8_1_MF8_3_MXS2_Mux4_1(in4087, M8_MF8_1_MF8_3_MXS2_Not_ContHi);
and3 M8_MF8_1_MF8_3_MXS2_Mux4_2(FXbus_7, M8_MF8_1_MF8_3_MXS2_Not_ContHi, M8_MF8_1_MF8_3_MXS2_Not_ContLo, M8_MF8_1_MF8_3_MXS2_line2);
and3 M8_MF8_1_MF8_3_MXS2_Mux4_3(FYbus_7, M8_MF8_1_MF8_3_MXS2_Not_ContHi, in4088, M8_MF8_1_MF8_3_MXS2_line3);
and3 M8_MF8_1_MF8_3_MXS2_Mux4_4(in46, in4087, M8_MF8_1_MF8_3_MXS2_Not_ContLo, M8_MF8_1_MF8_3_MXS2_line4);
and3 M8_MF8_1_MF8_3_MXS2_Mux4_5(in49, in4087, in4088, M8_MF8_1_MF8_3_MXS2_line5);
or4 M8_MF8_1_MF8_3_MXS2_Mux4_6(M8_MF8_1_MF8_3_MXS2_line2, M8_MF8_1_MF8_3_MXS2_line3, M8_MF8_1_MF8_3_MXS2_line4, M8_MF8_1_MF8_3_MXS2_line5, out732);
inv M8_MF8_1_MF8_3_MXS3_Mux4_0(in4089, M8_MF8_1_MF8_3_MXS3_Not_ContLo);
inv M8_MF8_1_MF8_3_MXS3_Mux4_1(in4090, M8_MF8_1_MF8_3_MXS3_Not_ContHi);
and3 M8_MF8_1_MF8_3_MXS3_Mux4_2(FXbus_7, M8_MF8_1_MF8_3_MXS3_Not_ContHi, M8_MF8_1_MF8_3_MXS3_Not_ContLo, M8_MF8_1_MF8_3_MXS3_line2);
and3 M8_MF8_1_MF8_3_MXS3_Mux4_3(FYbus_7, M8_MF8_1_MF8_3_MXS3_Not_ContHi, in4089, M8_MF8_1_MF8_3_MXS3_line3);
and3 M8_MF8_1_MF8_3_MXS3_Mux4_4(in46, in4090, M8_MF8_1_MF8_3_MXS3_Not_ContLo, M8_MF8_1_MF8_3_MXS3_line4);
and3 M8_MF8_1_MF8_3_MXS3_Mux4_5(in49, in4090, in4089, M8_MF8_1_MF8_3_MXS3_line5);
or4 M8_MF8_1_MF8_3_MXS3_Mux4_6(M8_MF8_1_MF8_3_MXS3_line2, M8_MF8_1_MF8_3_MXS3_line3, M8_MF8_1_MF8_3_MXS3_line4, M8_MF8_1_MF8_3_MXS3_line5, out772);
and2 M8_MF8_1_MF8_3_MXS4(M8_MF8_1_MF8_3_tempOut1, in137, out651);
and2 M8_MF8_1_MF8_3_MXS5(M8_MF8_1_MF8_3_tempOut2, in137, out685);
inv M8_MF8_2_MXS0_Mux4_0(in1689, M8_MF8_2_MXS0_Not_ContLo);
inv M8_MF8_2_MXS0_Mux4_1(in1690, M8_MF8_2_MXS0_Not_ContHi);
and3 M8_MF8_2_MXS0_Mux4_2(FXbus_8, M8_MF8_2_MXS0_Not_ContHi, M8_MF8_2_MXS0_Not_ContLo, M8_MF8_2_MXS0_line2);
and3 M8_MF8_2_MXS0_Mux4_3(FYbus_8, M8_MF8_2_MXS0_Not_ContHi, in1689, M8_MF8_2_MXS0_line3);
and3 M8_MF8_2_MXS0_Mux4_4(in191, in1690, M8_MF8_2_MXS0_Not_ContLo, M8_MF8_2_MXS0_line4);
and3 M8_MF8_2_MXS0_Mux4_5(in161, in1690, in1689, M8_MF8_2_MXS0_line5);
or4 M8_MF8_2_MXS0_Mux4_6(M8_MF8_2_MXS0_line2, M8_MF8_2_MXS0_line3, M8_MF8_2_MXS0_line4, M8_MF8_2_MXS0_line5, M8_MF8_2_tempOut1);
inv M8_MF8_2_MXS1_Mux4_0(in1691, M8_MF8_2_MXS1_Not_ContLo);
inv M8_MF8_2_MXS1_Mux4_1(in1694, M8_MF8_2_MXS1_Not_ContHi);
and3 M8_MF8_2_MXS1_Mux4_2(FXbus_8, M8_MF8_2_MXS1_Not_ContHi, M8_MF8_2_MXS1_Not_ContLo, M8_MF8_2_MXS1_line2);
and3 M8_MF8_2_MXS1_Mux4_3(FYbus_8, M8_MF8_2_MXS1_Not_ContHi, in1691, M8_MF8_2_MXS1_line3);
and3 M8_MF8_2_MXS1_Mux4_4(in191, in1694, M8_MF8_2_MXS1_Not_ContLo, M8_MF8_2_MXS1_line4);
and3 M8_MF8_2_MXS1_Mux4_5(in161, in1694, in1691, M8_MF8_2_MXS1_line5);
or4 M8_MF8_2_MXS1_Mux4_6(M8_MF8_2_MXS1_line2, M8_MF8_2_MXS1_line3, M8_MF8_2_MXS1_line4, M8_MF8_2_MXS1_line5, M8_MF8_2_tempOut2);
inv M8_MF8_2_MXS2_Mux4_0(in4088, M8_MF8_2_MXS2_Not_ContLo);
inv M8_MF8_2_MXS2_Mux4_1(in4087, M8_MF8_2_MXS2_Not_ContHi);
and3 M8_MF8_2_MXS2_Mux4_2(FXbus_8, M8_MF8_2_MXS2_Not_ContHi, M8_MF8_2_MXS2_Not_ContLo, M8_MF8_2_MXS2_line2);
and3 M8_MF8_2_MXS2_Mux4_3(FYbus_8, M8_MF8_2_MXS2_Not_ContHi, in4088, M8_MF8_2_MXS2_line3);
and3 M8_MF8_2_MXS2_Mux4_4(in109, in4087, M8_MF8_2_MXS2_Not_ContLo, M8_MF8_2_MXS2_line4);
and3 M8_MF8_2_MXS2_Mux4_5(in106, in4087, in4088, M8_MF8_2_MXS2_line5);
or4 M8_MF8_2_MXS2_Mux4_6(M8_MF8_2_MXS2_line2, M8_MF8_2_MXS2_line3, M8_MF8_2_MXS2_line4, M8_MF8_2_MXS2_line5, out727);
inv M8_MF8_2_MXS3_Mux4_0(in4089, M8_MF8_2_MXS3_Not_ContLo);
inv M8_MF8_2_MXS3_Mux4_1(in4090, M8_MF8_2_MXS3_Not_ContHi);
and3 M8_MF8_2_MXS3_Mux4_2(FXbus_8, M8_MF8_2_MXS3_Not_ContHi, M8_MF8_2_MXS3_Not_ContLo, M8_MF8_2_MXS3_line2);
and3 M8_MF8_2_MXS3_Mux4_3(FYbus_8, M8_MF8_2_MXS3_Not_ContHi, in4089, M8_MF8_2_MXS3_line3);
and3 M8_MF8_2_MXS3_Mux4_4(in109, in4090, M8_MF8_2_MXS3_Not_ContLo, M8_MF8_2_MXS3_line4);
and3 M8_MF8_2_MXS3_Mux4_5(in106, in4090, in4089, M8_MF8_2_MXS3_line5);
or4 M8_MF8_2_MXS3_Mux4_6(M8_MF8_2_MXS3_line2, M8_MF8_2_MXS3_line3, M8_MF8_2_MXS3_line4, M8_MF8_2_MXS3_line5, out712);
and2 M8_MF8_2_MXS4(M8_MF8_2_tempOut1, in137, out654);
and2 M8_MF8_2_MXS5(M8_MF8_2_tempOut2, in137, out688);
inv M9_Inv9_0_Inv4_0(FXbus_0, out822);
inv M9_Inv9_0_Inv4_1(FXbus_1, out838);
inv M9_Inv9_0_Inv4_2(FXbus_2, out836);
inv M9_Inv9_0_Inv4_3(FXbus_3, out834);
inv M9_Inv9_1_Inv4_0(FXbus_4, out832);
inv M9_Inv9_1_Inv4_1(FXbus_5, out830);
inv M9_Inv9_1_Inv4_2(FXbus_6, out828);
inv M9_Inv9_1_Inv4_3(FXbus_7, out826);
inv M9_Inv9_2(FXbus_8, out824);
inv M10_Inv9_0_Inv4_0(FYbus_0, out861);
inv M10_Inv9_0_Inv4_1(FYbus_1, out877);
inv M10_Inv9_0_Inv4_2(FYbus_2, out875);
inv M10_Inv9_0_Inv4_3(FYbus_3, out873);
inv M10_Inv9_1_Inv4_0(FYbus_4, out871);
inv M10_Inv9_1_Inv4_1(FYbus_5, out869);
inv M10_Inv9_1_Inv4_2(FYbus_6, out867);
inv M10_Inv9_1_Inv4_3(FYbus_7, out865);
inv M10_Inv9_2(FYbus_8, out863);
nor9 M11_ZF0_n9(SumXbus_0, SumXbus_1, SumXbus_2, SumXbus_3, SumXbus_4, SumXbus_5, SumXbus_6, SumXbus_7, SumXbus_8, out585);
nor9 M11_ZF1_n9(SumYbus_0, SumYbus_1, SumYbus_2, SumYbus_3, SumYbus_4, SumYbus_5, SumYbus_6, SumYbus_7, SumYbus_8, out575);
nor9 M11_ZF2_n9(LogicXbus_0, LogicXbus_1, LogicXbus_2, LogicXbus_3, LogicXbus_4, LogicXbus_5, LogicXbus_6, LogicXbus_7, LogicXbus_8, out598);
nor9 M11_ZF3_n9(LogicYbus_0, LogicYbus_1, LogicYbus_2, LogicYbus_3, LogicYbus_4, LogicYbus_5, LogicYbus_6, LogicYbus_7, LogicYbus_8, out610);
inv M12_BPC0_Mux2_0(in332, M12_BPC0_Not_ContIn);
and2 M12_BPC0_Mux2_1(in369, M12_BPC0_Not_ContIn, M12_BPC0_line1);
and2 M12_BPC0_Mux2_2(in372, in332, M12_BPC0_line2);
or2 M12_BPC0_Mux2_3(M12_BPC0_line1, M12_BPC0_line2, M12_ParX);
inv M12_BPC1_Mux2_0(in335, M12_BPC1_Not_ContIn);
and2 M12_BPC1_Mux2_1(in289, M12_BPC1_Not_ContIn, M12_BPC1_line1);
and2 M12_BPC1_Mux2_2(in292, in335, M12_BPC1_line2);
or2 M12_BPC1_Mux2_3(M12_BPC1_line1, M12_BPC1_line2, M12_ParY);
inv M12_BPC2_PT0_Xo0(Xbus_5, M12_BPC2_PT0_NotA);
inv M12_BPC2_PT0_Xo1(Xbus_6, M12_BPC2_PT0_NotB);
nand2 M12_BPC2_PT0_Xo2(M12_BPC2_PT0_NotA, Xbus_6, M12_BPC2_PT0_line2);
nand2 M12_BPC2_PT0_Xo3(M12_BPC2_PT0_NotB, Xbus_5, M12_BPC2_PT0_line3);
nand2 M12_BPC2_PT0_Xo4(M12_BPC2_PT0_line2, M12_BPC2_PT0_line3, M12_BPC2_line0);
inv M12_BPC2_PT1_Xo0(Xbus_7, M12_BPC2_PT1_NotA);
inv M12_BPC2_PT1_Xo1(Xbus_8, M12_BPC2_PT1_NotB);
nand2 M12_BPC2_PT1_Xo2(M12_BPC2_PT1_NotA, Xbus_8, M12_BPC2_PT1_line2);
nand2 M12_BPC2_PT1_Xo3(M12_BPC2_PT1_NotB, Xbus_7, M12_BPC2_PT1_line3);
nand2 M12_BPC2_PT1_Xo4(M12_BPC2_PT1_line2, M12_BPC2_PT1_line3, M12_BPC2_line1);
inv M12_BPC2_PT2_Xo0(Xbus_0, M12_BPC2_PT2_NotA);
inv M12_BPC2_PT2_Xo1(M12_ParX, M12_BPC2_PT2_NotB);
nand2 M12_BPC2_PT2_Xo2(M12_BPC2_PT2_NotA, M12_ParX, M12_BPC2_PT2_line2);
nand2 M12_BPC2_PT2_Xo3(M12_BPC2_PT2_NotB, Xbus_0, M12_BPC2_PT2_line3);
nand2 M12_BPC2_PT2_Xo4(M12_BPC2_PT2_line2, M12_BPC2_PT2_line3, M12_BPC2_line2);
inv M12_BPC2_PT3_Xo0(Xbus_1, M12_BPC2_PT3_NotA);
inv M12_BPC2_PT3_Xo1(Xbus_2, M12_BPC2_PT3_NotB);
nand2 M12_BPC2_PT3_Xo2(M12_BPC2_PT3_NotA, Xbus_2, M12_BPC2_PT3_line2);
nand2 M12_BPC2_PT3_Xo3(M12_BPC2_PT3_NotB, Xbus_1, M12_BPC2_PT3_line3);
nand2 M12_BPC2_PT3_Xo4(M12_BPC2_PT3_line2, M12_BPC2_PT3_line3, M12_BPC2_line3);
inv M12_BPC2_PT4_Xo0(Xbus_3, M12_BPC2_PT4_NotA);
inv M12_BPC2_PT4_Xo1(Xbus_4, M12_BPC2_PT4_NotB);
nand2 M12_BPC2_PT4_Xo2(M12_BPC2_PT4_NotA, Xbus_4, M12_BPC2_PT4_line2);
nand2 M12_BPC2_PT4_Xo3(M12_BPC2_PT4_NotB, Xbus_3, M12_BPC2_PT4_line3);
nand2 M12_BPC2_PT4_Xo4(M12_BPC2_PT4_line2, M12_BPC2_PT4_line3, M12_BPC2_line4);
inv M12_BPC2_PT5_Xo0(M12_BPC2_line0, M12_BPC2_PT5_NotA);
inv M12_BPC2_PT5_Xo1(M12_BPC2_line1, M12_BPC2_PT5_NotB);
nand2 M12_BPC2_PT5_Xo2(M12_BPC2_PT5_NotA, M12_BPC2_line1, M12_BPC2_PT5_line2);
nand2 M12_BPC2_PT5_Xo3(M12_BPC2_PT5_NotB, M12_BPC2_line0, M12_BPC2_PT5_line3);
nand2 M12_BPC2_PT5_Xo4(M12_BPC2_PT5_line2, M12_BPC2_PT5_line3, M12_BPC2_line5);
inv M12_BPC2_PT6_Xo3_0(M12_BPC2_line2, M12_BPC2_PT6_NotA);
inv M12_BPC2_PT6_Xo3_1(M12_BPC2_line3, M12_BPC2_PT6_NotB);
inv M12_BPC2_PT6_Xo3_2(M12_BPC2_line4, M12_BPC2_PT6_NotC);
and3 M12_BPC2_PT6_Xo3_3(M12_BPC2_PT6_NotA, M12_BPC2_PT6_NotB, M12_BPC2_line4, M12_BPC2_PT6_line3);
and3 M12_BPC2_PT6_Xo3_4(M12_BPC2_PT6_NotA, M12_BPC2_line3, M12_BPC2_PT6_NotC, M12_BPC2_PT6_line4);
and3 M12_BPC2_PT6_Xo3_5(M12_BPC2_line2, M12_BPC2_PT6_NotB, M12_BPC2_PT6_NotC, M12_BPC2_PT6_line5);
and3 M12_BPC2_PT6_Xo3_6(M12_BPC2_line2, M12_BPC2_line3, M12_BPC2_line4, M12_BPC2_PT6_line6);
nor2 M12_BPC2_PT6_Xo3_7(M12_BPC2_PT6_line3, M12_BPC2_PT6_line4, M12_BPC2_PT6_line7);
nor2 M12_BPC2_PT6_Xo3_8(M12_BPC2_PT6_line5, M12_BPC2_PT6_line6, M12_BPC2_PT6_line8);
nand2 M12_BPC2_PT6_Xo3_9(M12_BPC2_PT6_line7, M12_BPC2_PT6_line8, M12_BPC2_line6);
inv M12_BPC2_PT7_Xo0(M12_BPC2_line5, M12_BPC2_PT7_NotA);
inv M12_BPC2_PT7_Xo1(M12_BPC2_line6, M12_BPC2_PT7_NotB);
nand2 M12_BPC2_PT7_Xo2(M12_BPC2_PT7_NotA, M12_BPC2_line6, M12_BPC2_PT7_line2);
nand2 M12_BPC2_PT7_Xo3(M12_BPC2_PT7_NotB, M12_BPC2_line5, M12_BPC2_PT7_line3);
nand2 M12_BPC2_PT7_Xo4(M12_BPC2_PT7_line2, M12_BPC2_PT7_line3, out998);
inv M12_BPC3_PT0_Xo0(in316, M12_BPC3_PT0_NotA);
inv M12_BPC3_PT0_Xo1(in308, M12_BPC3_PT0_NotB);
nand2 M12_BPC3_PT0_Xo2(M12_BPC3_PT0_NotA, in308, M12_BPC3_PT0_line2);
nand2 M12_BPC3_PT0_Xo3(M12_BPC3_PT0_NotB, in316, M12_BPC3_PT0_line3);
nand2 M12_BPC3_PT0_Xo4(M12_BPC3_PT0_line2, M12_BPC3_PT0_line3, M12_BPC3_line0);
inv M12_BPC3_PT1_Xo0(in302, M12_BPC3_PT1_NotA);
inv M12_BPC3_PT1_Xo1(in293, M12_BPC3_PT1_NotB);
nand2 M12_BPC3_PT1_Xo2(M12_BPC3_PT1_NotA, in293, M12_BPC3_PT1_line2);
nand2 M12_BPC3_PT1_Xo3(M12_BPC3_PT1_NotB, in302, M12_BPC3_PT1_line3);
nand2 M12_BPC3_PT1_Xo4(M12_BPC3_PT1_line2, M12_BPC3_PT1_line3, M12_BPC3_line1);
inv M12_BPC3_PT2_Xo0(in361, M12_BPC3_PT2_NotA);
inv M12_BPC3_PT2_Xo1(in369, M12_BPC3_PT2_NotB);
nand2 M12_BPC3_PT2_Xo2(M12_BPC3_PT2_NotA, in369, M12_BPC3_PT2_line2);
nand2 M12_BPC3_PT2_Xo3(M12_BPC3_PT2_NotB, in361, M12_BPC3_PT2_line3);
nand2 M12_BPC3_PT2_Xo4(M12_BPC3_PT2_line2, M12_BPC3_PT2_line3, M12_BPC3_line2);
inv M12_BPC3_PT3_Xo0(in351, M12_BPC3_PT3_NotA);
inv M12_BPC3_PT3_Xo1(in341, M12_BPC3_PT3_NotB);
nand2 M12_BPC3_PT3_Xo2(M12_BPC3_PT3_NotA, in341, M12_BPC3_PT3_line2);
nand2 M12_BPC3_PT3_Xo3(M12_BPC3_PT3_NotB, in351, M12_BPC3_PT3_line3);
nand2 M12_BPC3_PT3_Xo4(M12_BPC3_PT3_line2, M12_BPC3_PT3_line3, M12_BPC3_line3);
inv M12_BPC3_PT4_Xo0(vdd, M12_BPC3_PT4_NotA);
inv M12_BPC3_PT4_Xo1(in324, M12_BPC3_PT4_NotB);
nand2 M12_BPC3_PT4_Xo2(M12_BPC3_PT4_NotA, in324, M12_BPC3_PT4_line2);
nand2 M12_BPC3_PT4_Xo3(M12_BPC3_PT4_NotB, vdd, M12_BPC3_PT4_line3);
nand2 M12_BPC3_PT4_Xo4(M12_BPC3_PT4_line2, M12_BPC3_PT4_line3, M12_BPC3_line4);
inv M12_BPC3_PT5_Xo0(M12_BPC3_line0, M12_BPC3_PT5_NotA);
inv M12_BPC3_PT5_Xo1(M12_BPC3_line1, M12_BPC3_PT5_NotB);
nand2 M12_BPC3_PT5_Xo2(M12_BPC3_PT5_NotA, M12_BPC3_line1, M12_BPC3_PT5_line2);
nand2 M12_BPC3_PT5_Xo3(M12_BPC3_PT5_NotB, M12_BPC3_line0, M12_BPC3_PT5_line3);
nand2 M12_BPC3_PT5_Xo4(M12_BPC3_PT5_line2, M12_BPC3_PT5_line3, M12_BPC3_line5);
inv M12_BPC3_PT6_Xo3_0(M12_BPC3_line2, M12_BPC3_PT6_NotA);
inv M12_BPC3_PT6_Xo3_1(M12_BPC3_line3, M12_BPC3_PT6_NotB);
inv M12_BPC3_PT6_Xo3_2(M12_BPC3_line4, M12_BPC3_PT6_NotC);
and3 M12_BPC3_PT6_Xo3_3(M12_BPC3_PT6_NotA, M12_BPC3_PT6_NotB, M12_BPC3_line4, M12_BPC3_PT6_line3);
and3 M12_BPC3_PT6_Xo3_4(M12_BPC3_PT6_NotA, M12_BPC3_line3, M12_BPC3_PT6_NotC, M12_BPC3_PT6_line4);
and3 M12_BPC3_PT6_Xo3_5(M12_BPC3_line2, M12_BPC3_PT6_NotB, M12_BPC3_PT6_NotC, M12_BPC3_PT6_line5);
and3 M12_BPC3_PT6_Xo3_6(M12_BPC3_line2, M12_BPC3_line3, M12_BPC3_line4, M12_BPC3_PT6_line6);
nor2 M12_BPC3_PT6_Xo3_7(M12_BPC3_PT6_line3, M12_BPC3_PT6_line4, M12_BPC3_PT6_line7);
nor2 M12_BPC3_PT6_Xo3_8(M12_BPC3_PT6_line5, M12_BPC3_PT6_line6, M12_BPC3_PT6_line8);
nand2 M12_BPC3_PT6_Xo3_9(M12_BPC3_PT6_line7, M12_BPC3_PT6_line8, M12_BPC3_line6);
inv M12_BPC3_PT7_Xo0(M12_BPC3_line5, M12_BPC3_PT7_NotA);
inv M12_BPC3_PT7_Xo1(M12_BPC3_line6, M12_BPC3_PT7_NotB);
nand2 M12_BPC3_PT7_Xo2(M12_BPC3_PT7_NotA, M12_BPC3_line6, M12_BPC3_PT7_line2);
nand2 M12_BPC3_PT7_Xo3(M12_BPC3_PT7_NotB, M12_BPC3_line5, M12_BPC3_PT7_line3);
nand2 M12_BPC3_PT7_Xo4(M12_BPC3_PT7_line2, M12_BPC3_PT7_line3, out1002);
inv M12_BPC4_PT0_Xo0(Ybus_5, M12_BPC4_PT0_NotA);
inv M12_BPC4_PT0_Xo1(Ybus_6, M12_BPC4_PT0_NotB);
nand2 M12_BPC4_PT0_Xo2(M12_BPC4_PT0_NotA, Ybus_6, M12_BPC4_PT0_line2);
nand2 M12_BPC4_PT0_Xo3(M12_BPC4_PT0_NotB, Ybus_5, M12_BPC4_PT0_line3);
nand2 M12_BPC4_PT0_Xo4(M12_BPC4_PT0_line2, M12_BPC4_PT0_line3, M12_BPC4_line0);
inv M12_BPC4_PT1_Xo0(Ybus_7, M12_BPC4_PT1_NotA);
inv M12_BPC4_PT1_Xo1(Ybus_8, M12_BPC4_PT1_NotB);
nand2 M12_BPC4_PT1_Xo2(M12_BPC4_PT1_NotA, Ybus_8, M12_BPC4_PT1_line2);
nand2 M12_BPC4_PT1_Xo3(M12_BPC4_PT1_NotB, Ybus_7, M12_BPC4_PT1_line3);
nand2 M12_BPC4_PT1_Xo4(M12_BPC4_PT1_line2, M12_BPC4_PT1_line3, M12_BPC4_line1);
inv M12_BPC4_PT2_Xo0(Ybus_0, M12_BPC4_PT2_NotA);
inv M12_BPC4_PT2_Xo1(M12_ParY, M12_BPC4_PT2_NotB);
nand2 M12_BPC4_PT2_Xo2(M12_BPC4_PT2_NotA, M12_ParY, M12_BPC4_PT2_line2);
nand2 M12_BPC4_PT2_Xo3(M12_BPC4_PT2_NotB, Ybus_0, M12_BPC4_PT2_line3);
nand2 M12_BPC4_PT2_Xo4(M12_BPC4_PT2_line2, M12_BPC4_PT2_line3, M12_BPC4_line2);
inv M12_BPC4_PT3_Xo0(Ybus_1, M12_BPC4_PT3_NotA);
inv M12_BPC4_PT3_Xo1(Ybus_2, M12_BPC4_PT3_NotB);
nand2 M12_BPC4_PT3_Xo2(M12_BPC4_PT3_NotA, Ybus_2, M12_BPC4_PT3_line2);
nand2 M12_BPC4_PT3_Xo3(M12_BPC4_PT3_NotB, Ybus_1, M12_BPC4_PT3_line3);
nand2 M12_BPC4_PT3_Xo4(M12_BPC4_PT3_line2, M12_BPC4_PT3_line3, M12_BPC4_line3);
inv M12_BPC4_PT4_Xo0(Ybus_3, M12_BPC4_PT4_NotA);
inv M12_BPC4_PT4_Xo1(Ybus_4, M12_BPC4_PT4_NotB);
nand2 M12_BPC4_PT4_Xo2(M12_BPC4_PT4_NotA, Ybus_4, M12_BPC4_PT4_line2);
nand2 M12_BPC4_PT4_Xo3(M12_BPC4_PT4_NotB, Ybus_3, M12_BPC4_PT4_line3);
nand2 M12_BPC4_PT4_Xo4(M12_BPC4_PT4_line2, M12_BPC4_PT4_line3, M12_BPC4_line4);
inv M12_BPC4_PT5_Xo0(M12_BPC4_line0, M12_BPC4_PT5_NotA);
inv M12_BPC4_PT5_Xo1(M12_BPC4_line1, M12_BPC4_PT5_NotB);
nand2 M12_BPC4_PT5_Xo2(M12_BPC4_PT5_NotA, M12_BPC4_line1, M12_BPC4_PT5_line2);
nand2 M12_BPC4_PT5_Xo3(M12_BPC4_PT5_NotB, M12_BPC4_line0, M12_BPC4_PT5_line3);
nand2 M12_BPC4_PT5_Xo4(M12_BPC4_PT5_line2, M12_BPC4_PT5_line3, M12_BPC4_line5);
inv M12_BPC4_PT6_Xo3_0(M12_BPC4_line2, M12_BPC4_PT6_NotA);
inv M12_BPC4_PT6_Xo3_1(M12_BPC4_line3, M12_BPC4_PT6_NotB);
inv M12_BPC4_PT6_Xo3_2(M12_BPC4_line4, M12_BPC4_PT6_NotC);
and3 M12_BPC4_PT6_Xo3_3(M12_BPC4_PT6_NotA, M12_BPC4_PT6_NotB, M12_BPC4_line4, M12_BPC4_PT6_line3);
and3 M12_BPC4_PT6_Xo3_4(M12_BPC4_PT6_NotA, M12_BPC4_line3, M12_BPC4_PT6_NotC, M12_BPC4_PT6_line4);
and3 M12_BPC4_PT6_Xo3_5(M12_BPC4_line2, M12_BPC4_PT6_NotB, M12_BPC4_PT6_NotC, M12_BPC4_PT6_line5);
and3 M12_BPC4_PT6_Xo3_6(M12_BPC4_line2, M12_BPC4_line3, M12_BPC4_line4, M12_BPC4_PT6_line6);
nor2 M12_BPC4_PT6_Xo3_7(M12_BPC4_PT6_line3, M12_BPC4_PT6_line4, M12_BPC4_PT6_line7);
nor2 M12_BPC4_PT6_Xo3_8(M12_BPC4_PT6_line5, M12_BPC4_PT6_line6, M12_BPC4_PT6_line8);
nand2 M12_BPC4_PT6_Xo3_9(M12_BPC4_PT6_line7, M12_BPC4_PT6_line8, M12_BPC4_line6);
inv M12_BPC4_PT7_Xo0(M12_BPC4_line5, M12_BPC4_PT7_NotA);
inv M12_BPC4_PT7_Xo1(M12_BPC4_line6, M12_BPC4_PT7_NotB);
nand2 M12_BPC4_PT7_Xo2(M12_BPC4_PT7_NotA, M12_BPC4_line6, M12_BPC4_PT7_line2);
nand2 M12_BPC4_PT7_Xo3(M12_BPC4_PT7_NotB, M12_BPC4_line5, M12_BPC4_PT7_line3);
nand2 M12_BPC4_PT7_Xo4(M12_BPC4_PT7_line2, M12_BPC4_PT7_line3, out1000);
inv M12_BPC5_PT0_Xo0(in226, M12_BPC5_PT0_NotA);
inv M12_BPC5_PT0_Xo1(in218, M12_BPC5_PT0_NotB);
nand2 M12_BPC5_PT0_Xo2(M12_BPC5_PT0_NotA, in218, M12_BPC5_PT0_line2);
nand2 M12_BPC5_PT0_Xo3(M12_BPC5_PT0_NotB, in226, M12_BPC5_PT0_line3);
nand2 M12_BPC5_PT0_Xo4(M12_BPC5_PT0_line2, M12_BPC5_PT0_line3, M12_BPC5_line0);
inv M12_BPC5_PT1_Xo0(in210, M12_BPC5_PT1_NotA);
inv M12_BPC5_PT1_Xo1(in206, M12_BPC5_PT1_NotB);
nand2 M12_BPC5_PT1_Xo2(M12_BPC5_PT1_NotA, in206, M12_BPC5_PT1_line2);
nand2 M12_BPC5_PT1_Xo3(M12_BPC5_PT1_NotB, in210, M12_BPC5_PT1_line3);
nand2 M12_BPC5_PT1_Xo4(M12_BPC5_PT1_line2, M12_BPC5_PT1_line3, M12_BPC5_line1);
inv M12_BPC5_PT2_Xo0(in281, M12_BPC5_PT2_NotA);
inv M12_BPC5_PT2_Xo1(in289, M12_BPC5_PT2_NotB);
nand2 M12_BPC5_PT2_Xo2(M12_BPC5_PT2_NotA, in289, M12_BPC5_PT2_line2);
nand2 M12_BPC5_PT2_Xo3(M12_BPC5_PT2_NotB, in281, M12_BPC5_PT2_line3);
nand2 M12_BPC5_PT2_Xo4(M12_BPC5_PT2_line2, M12_BPC5_PT2_line3, M12_BPC5_line2);
inv M12_BPC5_PT3_Xo0(in273, M12_BPC5_PT3_NotA);
inv M12_BPC5_PT3_Xo1(in265, M12_BPC5_PT3_NotB);
nand2 M12_BPC5_PT3_Xo2(M12_BPC5_PT3_NotA, in265, M12_BPC5_PT3_line2);
nand2 M12_BPC5_PT3_Xo3(M12_BPC5_PT3_NotB, in273, M12_BPC5_PT3_line3);
nand2 M12_BPC5_PT3_Xo4(M12_BPC5_PT3_line2, M12_BPC5_PT3_line3, M12_BPC5_line3);
inv M12_BPC5_PT4_Xo0(in257, M12_BPC5_PT4_NotA);
inv M12_BPC5_PT4_Xo1(in234, M12_BPC5_PT4_NotB);
nand2 M12_BPC5_PT4_Xo2(M12_BPC5_PT4_NotA, in234, M12_BPC5_PT4_line2);
nand2 M12_BPC5_PT4_Xo3(M12_BPC5_PT4_NotB, in257, M12_BPC5_PT4_line3);
nand2 M12_BPC5_PT4_Xo4(M12_BPC5_PT4_line2, M12_BPC5_PT4_line3, M12_BPC5_line4);
inv M12_BPC5_PT5_Xo0(M12_BPC5_line0, M12_BPC5_PT5_NotA);
inv M12_BPC5_PT5_Xo1(M12_BPC5_line1, M12_BPC5_PT5_NotB);
nand2 M12_BPC5_PT5_Xo2(M12_BPC5_PT5_NotA, M12_BPC5_line1, M12_BPC5_PT5_line2);
nand2 M12_BPC5_PT5_Xo3(M12_BPC5_PT5_NotB, M12_BPC5_line0, M12_BPC5_PT5_line3);
nand2 M12_BPC5_PT5_Xo4(M12_BPC5_PT5_line2, M12_BPC5_PT5_line3, M12_BPC5_line5);
inv M12_BPC5_PT6_Xo3_0(M12_BPC5_line2, M12_BPC5_PT6_NotA);
inv M12_BPC5_PT6_Xo3_1(M12_BPC5_line3, M12_BPC5_PT6_NotB);
inv M12_BPC5_PT6_Xo3_2(M12_BPC5_line4, M12_BPC5_PT6_NotC);
and3 M12_BPC5_PT6_Xo3_3(M12_BPC5_PT6_NotA, M12_BPC5_PT6_NotB, M12_BPC5_line4, M12_BPC5_PT6_line3);
and3 M12_BPC5_PT6_Xo3_4(M12_BPC5_PT6_NotA, M12_BPC5_line3, M12_BPC5_PT6_NotC, M12_BPC5_PT6_line4);
and3 M12_BPC5_PT6_Xo3_5(M12_BPC5_line2, M12_BPC5_PT6_NotB, M12_BPC5_PT6_NotC, M12_BPC5_PT6_line5);
and3 M12_BPC5_PT6_Xo3_6(M12_BPC5_line2, M12_BPC5_line3, M12_BPC5_line4, M12_BPC5_PT6_line6);
nor2 M12_BPC5_PT6_Xo3_7(M12_BPC5_PT6_line3, M12_BPC5_PT6_line4, M12_BPC5_PT6_line7);
nor2 M12_BPC5_PT6_Xo3_8(M12_BPC5_PT6_line5, M12_BPC5_PT6_line6, M12_BPC5_PT6_line8);
nand2 M12_BPC5_PT6_Xo3_9(M12_BPC5_PT6_line7, M12_BPC5_PT6_line8, M12_BPC5_line6);
inv M12_BPC5_PT7_Xo0(M12_BPC5_line5, M12_BPC5_PT7_NotA);
inv M12_BPC5_PT7_Xo1(M12_BPC5_line6, M12_BPC5_PT7_NotB);
nand2 M12_BPC5_PT7_Xo2(M12_BPC5_PT7_NotA, M12_BPC5_line6, M12_BPC5_PT7_line2);
nand2 M12_BPC5_PT7_Xo3(M12_BPC5_PT7_NotB, M12_BPC5_line5, M12_BPC5_PT7_line3);
nand2 M12_BPC5_PT7_Xo4(M12_BPC5_PT7_line2, M12_BPC5_PT7_line3, out1004);
inv M12_BPC6_Inv4_0(out1004, M12_NotParChk_0);
inv M12_BPC6_Inv4_1(out1000, M12_NotParChk_1);
inv M12_BPC6_Inv4_2(out1002, M12_NotParChk_2);
inv M12_BPC6_Inv4_3(out998, M12_NotParChk_3);
and5 M12_BPC7(M12_NotParChk_3, M12_NotParChk_2, M12_NotParChk_1, M12_NotParChk_0, in562, M12_line7);
and4 M12_BPC8(in386, in559, in556, in552, M12_line8);
and3 M12_BPC9(M12_line8, M12_line7, in245, out854);
and2 M13_UM13_0_MML0(in27, in31, M13_ContBeta);
inv M13_UM13_0_MML1(M13_ContBeta, M13_UM13_0_NotContBeta);
inv M13_UM13_0_MML2(in2358, M13_UM13_0_NotContIn2);
inv M13_UM13_0_MML3_Mux4_0_Mux2_0(M13_UM13_0_NotContIn2, M13_UM13_0_MML3_Mux4_0_Not_ContIn);
and2 M13_UM13_0_MML3_Mux4_0_Mux2_1(in34, M13_UM13_0_MML3_Mux4_0_Not_ContIn, M13_UM13_0_MML3_Mux4_0_line1);
and2 M13_UM13_0_MML3_Mux4_0_Mux2_2(in88, M13_UM13_0_NotContIn2, M13_UM13_0_MML3_Mux4_0_line2);
or2 M13_UM13_0_MML3_Mux4_0_Mux2_3(M13_UM13_0_MML3_Mux4_0_line1, M13_UM13_0_MML3_Mux4_0_line2, M13_UM13_0_tempOut1_0);
inv M13_UM13_0_MML3_Mux4_1_Mux2_0(M13_UM13_0_NotContIn2, M13_UM13_0_MML3_Mux4_1_Not_ContIn);
and2 M13_UM13_0_MML3_Mux4_1_Mux2_1(in34, M13_UM13_0_MML3_Mux4_1_Not_ContIn, M13_UM13_0_MML3_Mux4_1_line1);
and2 M13_UM13_0_MML3_Mux4_1_Mux2_2(in88, M13_UM13_0_NotContIn2, M13_UM13_0_MML3_Mux4_1_line2);
or2 M13_UM13_0_MML3_Mux4_1_Mux2_3(M13_UM13_0_MML3_Mux4_1_line1, M13_UM13_0_MML3_Mux4_1_line2, M13_UM13_0_tempOut1_1);
inv M13_UM13_0_MML3_Mux4_2_Mux2_0(M13_UM13_0_NotContIn2, M13_UM13_0_MML3_Mux4_2_Not_ContIn);
and2 M13_UM13_0_MML3_Mux4_2_Mux2_1(in83, M13_UM13_0_MML3_Mux4_2_Not_ContIn, M13_UM13_0_MML3_Mux4_2_line1);
and2 M13_UM13_0_MML3_Mux4_2_Mux2_2(in83, M13_UM13_0_NotContIn2, M13_UM13_0_MML3_Mux4_2_line2);
or2 M13_UM13_0_MML3_Mux4_2_Mux2_3(M13_UM13_0_MML3_Mux4_2_line1, M13_UM13_0_MML3_Mux4_2_line2, M13_UM13_0_tempOut1_2);
inv M13_UM13_0_MML3_Mux4_3_Mux2_0(M13_UM13_0_NotContIn2, M13_UM13_0_MML3_Mux4_3_Not_ContIn);
and2 M13_UM13_0_MML3_Mux4_3_Mux2_1(in87, M13_UM13_0_MML3_Mux4_3_Not_ContIn, M13_UM13_0_MML3_Mux4_3_line1);
and2 M13_UM13_0_MML3_Mux4_3_Mux2_2(in86, M13_UM13_0_NotContIn2, M13_UM13_0_MML3_Mux4_3_line2);
or2 M13_UM13_0_MML3_Mux4_3_Mux2_3(M13_UM13_0_MML3_Mux4_3_line1, M13_UM13_0_MML3_Mux4_3_line2, M13_UM13_0_tempOut1_3);
inv M13_UM13_0_MML4_Mx4_0_Mux4_0(in2358, M13_UM13_0_MML4_Mx4_0_Not_ContLo);
inv M13_UM13_0_MML4_Mx4_0_Mux4_1(M13_UM13_0_NotContBeta, M13_UM13_0_MML4_Mx4_0_Not_ContHi);
and3 M13_UM13_0_MML4_Mx4_0_Mux4_2(in26, M13_UM13_0_MML4_Mx4_0_Not_ContHi, M13_UM13_0_MML4_Mx4_0_Not_ContLo, M13_UM13_0_MML4_Mx4_0_line2);
and3 M13_UM13_0_MML4_Mx4_0_Mux4_3(in81, M13_UM13_0_MML4_Mx4_0_Not_ContHi, in2358, M13_UM13_0_MML4_Mx4_0_line3);
and3 M13_UM13_0_MML4_Mx4_0_Mux4_4(vdd, M13_UM13_0_NotContBeta, M13_UM13_0_MML4_Mx4_0_Not_ContLo, M13_UM13_0_MML4_Mx4_0_line4);
and3 M13_UM13_0_MML4_Mx4_0_Mux4_5(vdd, M13_UM13_0_NotContBeta, in2358, M13_UM13_0_MML4_Mx4_0_line5);
or4 M13_UM13_0_MML4_Mx4_0_Mux4_6(M13_UM13_0_MML4_Mx4_0_line2, M13_UM13_0_MML4_Mx4_0_line3, M13_UM13_0_MML4_Mx4_0_line4, M13_UM13_0_MML4_Mx4_0_line5, M13_UM13_0_tempOut2_0);
inv M13_UM13_0_MML4_Mx4_1_Mux4_0(in2358, M13_UM13_0_MML4_Mx4_1_Not_ContLo);
inv M13_UM13_0_MML4_Mx4_1_Mux4_1(M13_UM13_0_NotContBeta, M13_UM13_0_MML4_Mx4_1_Not_ContHi);
and3 M13_UM13_0_MML4_Mx4_1_Mux4_2(in24, M13_UM13_0_MML4_Mx4_1_Not_ContHi, M13_UM13_0_MML4_Mx4_1_Not_ContLo, M13_UM13_0_MML4_Mx4_1_line2);
and3 M13_UM13_0_MML4_Mx4_1_Mux4_3(in25, M13_UM13_0_MML4_Mx4_1_Not_ContHi, in2358, M13_UM13_0_MML4_Mx4_1_line3);
and3 M13_UM13_0_MML4_Mx4_1_Mux4_4(vdd, M13_UM13_0_NotContBeta, M13_UM13_0_MML4_Mx4_1_Not_ContLo, M13_UM13_0_MML4_Mx4_1_line4);
and3 M13_UM13_0_MML4_Mx4_1_Mux4_5(vdd, M13_UM13_0_NotContBeta, in2358, M13_UM13_0_MML4_Mx4_1_line5);
or4 M13_UM13_0_MML4_Mx4_1_Mux4_6(M13_UM13_0_MML4_Mx4_1_line2, M13_UM13_0_MML4_Mx4_1_line3, M13_UM13_0_MML4_Mx4_1_line4, M13_UM13_0_MML4_Mx4_1_line5, M13_UM13_0_tempOut2_1);
inv M13_UM13_0_MML4_Mx4_2_Mux4_0(in2358, M13_UM13_0_MML4_Mx4_2_Not_ContLo);
inv M13_UM13_0_MML4_Mx4_2_Mux4_1(M13_UM13_0_NotContBeta, M13_UM13_0_MML4_Mx4_2_Not_ContHi);
and3 M13_UM13_0_MML4_Mx4_2_Mux4_2(in82, M13_UM13_0_MML4_Mx4_2_Not_ContHi, M13_UM13_0_MML4_Mx4_2_Not_ContLo, M13_UM13_0_MML4_Mx4_2_line2);
and3 M13_UM13_0_MML4_Mx4_2_Mux4_3(in80, M13_UM13_0_MML4_Mx4_2_Not_ContHi, in2358, M13_UM13_0_MML4_Mx4_2_line3);
and3 M13_UM13_0_MML4_Mx4_2_Mux4_4(vdd, M13_UM13_0_NotContBeta, M13_UM13_0_MML4_Mx4_2_Not_ContLo, M13_UM13_0_MML4_Mx4_2_line4);
and3 M13_UM13_0_MML4_Mx4_2_Mux4_5(vdd, M13_UM13_0_NotContBeta, in2358, M13_UM13_0_MML4_Mx4_2_line5);
or4 M13_UM13_0_MML4_Mx4_2_Mux4_6(M13_UM13_0_MML4_Mx4_2_line2, M13_UM13_0_MML4_Mx4_2_line3, M13_UM13_0_MML4_Mx4_2_line4, M13_UM13_0_MML4_Mx4_2_line5, M13_UM13_0_tempOut2_2);
inv M13_UM13_0_MML4_Mx4_3_Mux4_0(in2358, M13_UM13_0_MML4_Mx4_3_Not_ContLo);
inv M13_UM13_0_MML4_Mx4_3_Mux4_1(M13_UM13_0_NotContBeta, M13_UM13_0_MML4_Mx4_3_Not_ContHi);
and3 M13_UM13_0_MML4_Mx4_3_Mux4_2(in79, M13_UM13_0_MML4_Mx4_3_Not_ContHi, M13_UM13_0_MML4_Mx4_3_Not_ContLo, M13_UM13_0_MML4_Mx4_3_line2);
and3 M13_UM13_0_MML4_Mx4_3_Mux4_3(in23, M13_UM13_0_MML4_Mx4_3_Not_ContHi, in2358, M13_UM13_0_MML4_Mx4_3_line3);
and3 M13_UM13_0_MML4_Mx4_3_Mux4_4(vdd, M13_UM13_0_NotContBeta, M13_UM13_0_MML4_Mx4_3_Not_ContLo, M13_UM13_0_MML4_Mx4_3_line4);
and3 M13_UM13_0_MML4_Mx4_3_Mux4_5(vdd, M13_UM13_0_NotContBeta, in2358, M13_UM13_0_MML4_Mx4_3_line5);
or4 M13_UM13_0_MML4_Mx4_3_Mux4_6(M13_UM13_0_MML4_Mx4_3_line2, M13_UM13_0_MML4_Mx4_3_line3, M13_UM13_0_MML4_Mx4_3_line4, M13_UM13_0_MML4_Mx4_3_line5, M13_UM13_0_tempOut2_3);
and2 M13_UM13_0_MML5_Ma0(M13_UM13_0_tempOut1_0, M13_ContBeta, M13_UM13_0_tempOut3_0);
and2 M13_UM13_0_MML5_Ma1(M13_UM13_0_tempOut1_1, M13_ContBeta, M13_UM13_0_tempOut3_1);
and2 M13_UM13_0_MML5_Ma2(M13_UM13_0_tempOut1_2, M13_ContBeta, M13_UM13_0_tempOut3_2);
and2 M13_UM13_0_MML5_Ma3(M13_UM13_0_tempOut1_3, M13_ContBeta, M13_UM13_0_tempOut3_3);
inv M13_UM13_0_MML6_Inv4_0(M13_UM13_0_tempOut3_0, out704);
inv M13_UM13_0_MML6_Inv4_1(M13_UM13_0_tempOut3_1, out717);
inv M13_UM13_0_MML6_Inv4_2(M13_UM13_0_tempOut3_2, out820);
inv M13_UM13_0_MML6_Inv4_3(M13_UM13_0_tempOut3_3, out636);
and2 M13_UM13_0_MML7_Ma0(M13_UM13_0_tempOut2_0, in141, out673);
and2 M13_UM13_0_MML7_Ma1(M13_UM13_0_tempOut2_1, in141, out639);
and2 M13_UM13_0_MML7_Ma2(M13_UM13_0_tempOut2_2, in141, out715);
and2 M13_UM13_0_MML7_Ma3(M13_UM13_0_tempOut2_3, in141, out707);
inv M13_UM13_0_MML8(Xbus_8, M13_UM13_0_NotMuxIn20);
nand2 M13_UM13_0_MML9_Xo0(M13_UM13_0_NotMuxIn20, in132, M13_UM13_0_MML9_NotAB);
and2 M13_UM13_0_MML9_Xo1(M13_UM13_0_NotMuxIn20, M13_UM13_0_MML9_NotAB, M13_UM13_0_MML9_line1);
and2 M13_UM13_0_MML9_Xo2(M13_UM13_0_MML9_NotAB, in132, M13_UM13_0_MML9_line2);
or2 M13_UM13_0_MML9_Xo3(M13_UM13_0_MML9_line1, M13_UM13_0_MML9_line2, M13_UM13_0_tempMuxin);
inv M13_UM13_0_MML10_Mux4_0(in3724, M13_UM13_0_MML10_Not_ContLo);
inv M13_UM13_0_MML10_Mux4_1(in3717, M13_UM13_0_MML10_Not_ContHi);
and3 M13_UM13_0_MML10_Mux4_2(LogicXbus_8, M13_UM13_0_MML10_Not_ContHi, M13_UM13_0_MML10_Not_ContLo, M13_UM13_0_MML10_line2);
and3 M13_UM13_0_MML10_Mux4_3(M13_UM13_0_tempMuxin, M13_UM13_0_MML10_Not_ContHi, in3724, M13_UM13_0_MML10_line3);
and3 M13_UM13_0_MML10_Mux4_4(in123, in3717, M13_UM13_0_MML10_Not_ContLo, M13_UM13_0_MML10_line4);
and3 M13_UM13_0_MML10_Mux4_5(SumXbus_8, in3717, in3724, M13_UM13_0_MML10_line5);
or4 M13_UM13_0_MML10_Mux4_6(M13_UM13_0_MML10_line2, M13_UM13_0_MML10_line3, M13_UM13_0_MML10_line4, M13_UM13_0_MML10_line5, M13_UM13_0_tempMuxout);
nand2 M13_UM13_0_MML11(in135, in4115, M13_UM13_0_tempMuxcont);
and2 M13_UM13_0_MML12(M13_UM13_0_tempMuxcont, M13_UM13_0_tempMuxout, out818);
nand2 M13_UM13_0_MML13_Xo0(M13_UM13_0_tempMuxin, SumXbus_8, M13_UM13_0_MML13_NotAB);
and2 M13_UM13_0_MML13_Xo1(M13_UM13_0_tempMuxin, M13_UM13_0_MML13_NotAB, M13_UM13_0_MML13_line1);
and2 M13_UM13_0_MML13_Xo2(M13_UM13_0_MML13_NotAB, SumXbus_8, M13_UM13_0_MML13_line2);
or2 M13_UM13_0_MML13_Xo3(M13_UM13_0_MML13_line1, M13_UM13_0_MML13_line2, out813);
inv M13_UM13_0_MML14(SumXbus_8, out623);
nand2 M13_UM13_1_MRL0(M13_ContBeta, in140, out656);
inv M13_UM13_1_MRL1(in2824, M13_UM13_1_NotMisc1);
and2 M13_UM13_1_MRL2(M13_UM13_1_NotMisc1, in27, M13_UM13_1_line2);
inv M13_UM13_1_MRL3(M13_UM13_1_line2, out845);
and2 M13_UM13_1_MRL4(in141, in145, out810);
nand2 M13_UM13_1_MRL5(in373, in1, M13_UM13_1_line6);
inv M13_UM13_1_MRL6(M13_UM13_1_line6, out634);
inv M13_UM13_1_MRL7(in3173, M13_UM13_1_NotMisc6);
and2 M13_UM13_1_MRL8(in136, M13_UM13_1_NotMisc6, out815);
and2 M13_UM13_1_MRL9(in386, in556, M13_UM13_1_line12);
inv M13_UM13_1_MRL10(M13_UM13_1_line12, out847);
and2 M13_UM13_1_MRL11(in552, in562, out601);
buffer M13_UM13_1_MRL12_B7_0(in141, out144);
buffer M13_UM13_1_MRL12_B7_1(in1, out993);
buffer M13_UM13_1_MRL12_B7_2(in3173, out973);
buffer M13_UM13_1_MRL12_B7_3(in549, out892);
buffer M13_UM13_1_MRL12_B7_4(in137, out926);
buffer M13_UM13_1_MRL12_B7_5(in293, out298);
buffer M13_UM13_1_MRL12_B7_6(in299, out887);
inv M13_UM13_1_MRL13_Inv4_0(in559, out851);
inv M13_UM13_1_MRL13_Inv4_1(in552, out849);
inv M13_UM13_1_MRL13_Inv4_2(in245, out848);
inv M13_UM13_1_MRL13_Inv4_3(in562, out850);
inv M13_UM13_1_MRL14_Inv4_0(in366, out600);
inv M13_UM13_1_MRL14_Inv4_1(in358, out612);
inv M13_UM13_1_MRL14_Inv4_2(in348, out599);
inv M13_UM13_1_MRL14_Inv4_3(in338, out611);
inv M13_UM13_1_MRL15_Inv4_0(M13_ContBeta, out809);
inv M13_UM13_1_MRL15_Inv4_1(in549, out602);
inv M13_UM13_1_MRL15_Inv4_2(in545, out594);
inv M13_UM13_1_MRL15_Inv4_3(in299, out593);

assign out618 = out629;
assign out621 = out591;
assign out626 = out615;
assign out632 = out588;
assign out923 = out144;
assign out939 = out993;
assign out921 = out993;
assign out978 = out993;
assign out949 = out993;
assign out889 = out887;
assign out603 = out594;
assign out604 = out594;
assign out606 = out602;
assign vdd = 1'b1;
assign gnd = 1'b0;

endmodule