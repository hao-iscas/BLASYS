module adder ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ,
    \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] ,
    \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] ,
    \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] ,
    \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] ,
    \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] ,
    \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] , \b[52] ,
    \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] , \b[60] ,
    \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] , \b[68] ,
    \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] , \b[76] ,
    \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] , \b[84] ,
    \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] ,
    \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127] , cOut  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] ,
    \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] ,
    \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] ,
    \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] ,
    \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] ,
    \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] ,
    \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] ,
    \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] ,
    \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] ,
    \b[68] , \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] ,
    \b[76] , \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] ,
    \b[84] , \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] ,
    \b[92] , \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] , cOut;
  wire n386, n387, n389, n390, n391, n392, n393, n394, n396, n397, n398,
    n399, n400, n401, n402, n404, n405, n406, n407, n408, n409, n410, n412,
    n413, n414, n415, n416, n417, n418, n420, n421, n422, n423, n424, n425,
    n426, n428, n429, n430, n431, n432, n433, n434, n436, n437, n438, n439,
    n440, n441, n442, n444, n445, n446, n447, n448, n449, n450, n452, n453,
    n454, n455, n456, n457, n458, n460, n461, n462, n463, n464, n465, n466,
    n468, n469, n470, n471, n472, n473, n474, n476, n477, n478, n479, n480,
    n481, n482, n484, n485, n486, n487, n488, n489, n490, n492, n493, n494,
    n495, n496, n497, n498, n500, n501, n502, n503, n504, n505, n506, n508,
    n509, n510, n511, n512, n513, n514, n516, n517, n518, n519, n520, n521,
    n522, n524, n525, n526, n527, n528, n529, n530, n532, n533, n534, n535,
    n536, n537, n538, n540, n541, n542, n543, n544, n545, n546, n548, n549,
    n550, n551, n552, n553, n554, n556, n557, n558, n559, n560, n561, n562,
    n564, n565, n566, n567, n568, n569, n570, n572, n573, n574, n575, n576,
    n577, n578, n580, n581, n582, n583, n584, n585, n586, n588, n589, n590,
    n591, n592, n593, n594, n596, n597, n598, n599, n600, n601, n602, n604,
    n605, n606, n607, n608, n609, n610, n612, n613, n614, n615, n616, n617,
    n618, n620, n621, n622, n623, n624, n625, n626, n628, n629, n630, n631,
    n632, n633, n634, n636, n637, n638, n639, n640, n641, n642, n644, n645,
    n646, n647, n648, n649, n650, n652, n653, n654, n655, n656, n657, n658,
    n660, n661, n662, n663, n664, n665, n666, n668, n669, n670, n671, n672,
    n673, n674, n676, n677, n678, n679, n680, n681, n682, n684, n685, n686,
    n687, n688, n689, n690, n692, n693, n694, n695, n696, n697, n698, n700,
    n701, n702, n703, n704, n705, n706, n708, n709, n710, n711, n712, n713,
    n714, n716, n717, n718, n719, n720, n721, n722, n724, n725, n726, n727,
    n728, n729, n730, n732, n733, n734, n735, n736, n737, n738, n740, n741,
    n742, n743, n744, n745, n746, n748, n749, n750, n751, n752, n753, n754,
    n756, n757, n758, n759, n760, n761, n762, n764, n765, n766, n767, n768,
    n769, n770, n772, n773, n774, n775, n776, n777, n778, n780, n781, n782,
    n783, n784, n785, n786, n788, n789, n790, n791, n792, n793, n794, n796,
    n797, n798, n799, n800, n801, n802, n804, n805, n806, n807, n808, n809,
    n810, n812, n813, n814, n815, n816, n817, n818, n820, n821, n822, n823,
    n824, n825, n826, n828, n829, n830, n831, n832, n833, n834, n836, n837,
    n838, n839, n840, n841, n842, n844, n845, n846, n847, n848, n849, n850,
    n852, n853, n854, n855, n856, n857, n858, n860, n861, n862, n863, n864,
    n865, n866, n868, n869, n870, n871, n872, n873, n874, n876, n877, n878,
    n879, n880, n881, n882, n884, n885, n886, n887, n888, n889, n890, n892,
    n893, n894, n895, n896, n897, n898, n900, n901, n902, n903, n904, n905,
    n906, n908, n909, n910, n911, n912, n913, n914, n916, n917, n918, n919,
    n920, n921, n922, n924, n925, n926, n927, n928, n929, n930, n932, n933,
    n934, n935, n936, n937, n938, n940, n941, n942, n943, n944, n945, n946,
    n948, n949, n950, n951, n952, n953, n954, n956, n957, n958, n959, n960,
    n961, n962, n964, n965, n966, n967, n968, n969, n970, n972, n973, n974,
    n975, n976, n977, n978, n980, n981, n982, n983, n984, n985, n986, n988,
    n989, n990, n991, n992, n993, n994, n996, n997, n998, n999, n1000,
    n1001, n1002, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1012,
    n1013, n1014, n1015, n1016, n1017, n1018, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
    n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1052, n1053, n1054, n1055, n1056, n1057,
    n1058, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098, n1100, n1101, n1102, n1103,
    n1104, n1105, n1106, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
    n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1172,
    n1173, n1174, n1175, n1176, n1177, n1178, n1180, n1181, n1182, n1183,
    n1184, n1185, n1186, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
    n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1204, n1205, n1206,
    n1207, n1208, n1209, n1210, n1212, n1213, n1214, n1215, n1216, n1217,
    n1218, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1236, n1237, n1238, n1239, n1240,
    n1241, n1242, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1252,
    n1253, n1254, n1255, n1256, n1257, n1258, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
    n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1292, n1293, n1294, n1295, n1296, n1297,
    n1298, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1316, n1317, n1318, n1319, n1320,
    n1321, n1322, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1332,
    n1333, n1334, n1335, n1336, n1337, n1338, n1340, n1341, n1342, n1343,
    n1344, n1345, n1346, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
    n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1364, n1365, n1366,
    n1367, n1368, n1369, n1370, n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1404;
  assign n386 = \a[0]  & ~\b[0] ;
  assign n387 = ~\a[0]  & \b[0] ;
  assign \f[0]  = n386 | n387;
  assign n389 = \a[0]  & \b[0] ;
  assign n390 = ~\a[1]  & ~\b[1] ;
  assign n391 = \a[1]  & \b[1] ;
  assign n392 = ~n390 & ~n391;
  assign n393 = n389 & ~n392;
  assign n394 = ~n389 & n392;
  assign \f[1]  = n393 | n394;
  assign n396 = n389 & ~n390;
  assign n397 = ~n391 & ~n396;
  assign n398 = ~\a[2]  & ~\b[2] ;
  assign n399 = \a[2]  & \b[2] ;
  assign n400 = ~n398 & ~n399;
  assign n401 = n397 & ~n400;
  assign n402 = ~n397 & n400;
  assign \f[2]  = ~n401 & ~n402;
  assign n404 = ~n397 & ~n398;
  assign n405 = ~n399 & ~n404;
  assign n406 = ~\a[3]  & ~\b[3] ;
  assign n407 = \a[3]  & \b[3] ;
  assign n408 = ~n406 & ~n407;
  assign n409 = n405 & ~n408;
  assign n410 = ~n405 & n408;
  assign \f[3]  = ~n409 & ~n410;
  assign n412 = ~n405 & ~n406;
  assign n413 = ~n407 & ~n412;
  assign n414 = ~\a[4]  & ~\b[4] ;
  assign n415 = \a[4]  & \b[4] ;
  assign n416 = ~n414 & ~n415;
  assign n417 = n413 & ~n416;
  assign n418 = ~n413 & n416;
  assign \f[4]  = ~n417 & ~n418;
  assign n420 = ~n413 & ~n414;
  assign n421 = ~n415 & ~n420;
  assign n422 = ~\a[5]  & ~\b[5] ;
  assign n423 = \a[5]  & \b[5] ;
  assign n424 = ~n422 & ~n423;
  assign n425 = n421 & ~n424;
  assign n426 = ~n421 & n424;
  assign \f[5]  = ~n425 & ~n426;
  assign n428 = ~n421 & ~n422;
  assign n429 = ~n423 & ~n428;
  assign n430 = ~\a[6]  & ~\b[6] ;
  assign n431 = \a[6]  & \b[6] ;
  assign n432 = ~n430 & ~n431;
  assign n433 = n429 & ~n432;
  assign n434 = ~n429 & n432;
  assign \f[6]  = ~n433 & ~n434;
  assign n436 = ~n429 & ~n430;
  assign n437 = ~n431 & ~n436;
  assign n438 = ~\a[7]  & ~\b[7] ;
  assign n439 = \a[7]  & \b[7] ;
  assign n440 = ~n438 & ~n439;
  assign n441 = n437 & ~n440;
  assign n442 = ~n437 & n440;
  assign \f[7]  = ~n441 & ~n442;
  assign n444 = ~n437 & ~n438;
  assign n445 = ~n439 & ~n444;
  assign n446 = ~\a[8]  & ~\b[8] ;
  assign n447 = \a[8]  & \b[8] ;
  assign n448 = ~n446 & ~n447;
  assign n449 = n445 & ~n448;
  assign n450 = ~n445 & n448;
  assign \f[8]  = ~n449 & ~n450;
  assign n452 = ~n445 & ~n446;
  assign n453 = ~n447 & ~n452;
  assign n454 = ~\a[9]  & ~\b[9] ;
  assign n455 = \a[9]  & \b[9] ;
  assign n456 = ~n454 & ~n455;
  assign n457 = n453 & ~n456;
  assign n458 = ~n453 & n456;
  assign \f[9]  = ~n457 & ~n458;
  assign n460 = ~n453 & ~n454;
  assign n461 = ~n455 & ~n460;
  assign n462 = ~\a[10]  & ~\b[10] ;
  assign n463 = \a[10]  & \b[10] ;
  assign n464 = ~n462 & ~n463;
  assign n465 = n461 & ~n464;
  assign n466 = ~n461 & n464;
  assign \f[10]  = ~n465 & ~n466;
  assign n468 = ~n461 & ~n462;
  assign n469 = ~n463 & ~n468;
  assign n470 = ~\a[11]  & ~\b[11] ;
  assign n471 = \a[11]  & \b[11] ;
  assign n472 = ~n470 & ~n471;
  assign n473 = n469 & ~n472;
  assign n474 = ~n469 & n472;
  assign \f[11]  = ~n473 & ~n474;
  assign n476 = ~n469 & ~n470;
  assign n477 = ~n471 & ~n476;
  assign n478 = ~\a[12]  & ~\b[12] ;
  assign n479 = \a[12]  & \b[12] ;
  assign n480 = ~n478 & ~n479;
  assign n481 = n477 & ~n480;
  assign n482 = ~n477 & n480;
  assign \f[12]  = ~n481 & ~n482;
  assign n484 = ~n477 & ~n478;
  assign n485 = ~n479 & ~n484;
  assign n486 = ~\a[13]  & ~\b[13] ;
  assign n487 = \a[13]  & \b[13] ;
  assign n488 = ~n486 & ~n487;
  assign n489 = n485 & ~n488;
  assign n490 = ~n485 & n488;
  assign \f[13]  = ~n489 & ~n490;
  assign n492 = ~n485 & ~n486;
  assign n493 = ~n487 & ~n492;
  assign n494 = ~\a[14]  & ~\b[14] ;
  assign n495 = \a[14]  & \b[14] ;
  assign n496 = ~n494 & ~n495;
  assign n497 = n493 & ~n496;
  assign n498 = ~n493 & n496;
  assign \f[14]  = ~n497 & ~n498;
  assign n500 = ~n493 & ~n494;
  assign n501 = ~n495 & ~n500;
  assign n502 = ~\a[15]  & ~\b[15] ;
  assign n503 = \a[15]  & \b[15] ;
  assign n504 = ~n502 & ~n503;
  assign n505 = n501 & ~n504;
  assign n506 = ~n501 & n504;
  assign \f[15]  = ~n505 & ~n506;
  assign n508 = ~n501 & ~n502;
  assign n509 = ~n503 & ~n508;
  assign n510 = ~\a[16]  & ~\b[16] ;
  assign n511 = \a[16]  & \b[16] ;
  assign n512 = ~n510 & ~n511;
  assign n513 = n509 & ~n512;
  assign n514 = ~n509 & n512;
  assign \f[16]  = ~n513 & ~n514;
  assign n516 = ~n509 & ~n510;
  assign n517 = ~n511 & ~n516;
  assign n518 = ~\a[17]  & ~\b[17] ;
  assign n519 = \a[17]  & \b[17] ;
  assign n520 = ~n518 & ~n519;
  assign n521 = n517 & ~n520;
  assign n522 = ~n517 & n520;
  assign \f[17]  = ~n521 & ~n522;
  assign n524 = ~n517 & ~n518;
  assign n525 = ~n519 & ~n524;
  assign n526 = ~\a[18]  & ~\b[18] ;
  assign n527 = \a[18]  & \b[18] ;
  assign n528 = ~n526 & ~n527;
  assign n529 = n525 & ~n528;
  assign n530 = ~n525 & n528;
  assign \f[18]  = ~n529 & ~n530;
  assign n532 = ~n525 & ~n526;
  assign n533 = ~n527 & ~n532;
  assign n534 = ~\a[19]  & ~\b[19] ;
  assign n535 = \a[19]  & \b[19] ;
  assign n536 = ~n534 & ~n535;
  assign n537 = n533 & ~n536;
  assign n538 = ~n533 & n536;
  assign \f[19]  = ~n537 & ~n538;
  assign n540 = ~n533 & ~n534;
  assign n541 = ~n535 & ~n540;
  assign n542 = ~\a[20]  & ~\b[20] ;
  assign n543 = \a[20]  & \b[20] ;
  assign n544 = ~n542 & ~n543;
  assign n545 = n541 & ~n544;
  assign n546 = ~n541 & n544;
  assign \f[20]  = ~n545 & ~n546;
  assign n548 = ~n541 & ~n542;
  assign n549 = ~n543 & ~n548;
  assign n550 = ~\a[21]  & ~\b[21] ;
  assign n551 = \a[21]  & \b[21] ;
  assign n552 = ~n550 & ~n551;
  assign n553 = n549 & ~n552;
  assign n554 = ~n549 & n552;
  assign \f[21]  = ~n553 & ~n554;
  assign n556 = ~n549 & ~n550;
  assign n557 = ~n551 & ~n556;
  assign n558 = ~\a[22]  & ~\b[22] ;
  assign n559 = \a[22]  & \b[22] ;
  assign n560 = ~n558 & ~n559;
  assign n561 = n557 & ~n560;
  assign n562 = ~n557 & n560;
  assign \f[22]  = ~n561 & ~n562;
  assign n564 = ~n557 & ~n558;
  assign n565 = ~n559 & ~n564;
  assign n566 = ~\a[23]  & ~\b[23] ;
  assign n567 = \a[23]  & \b[23] ;
  assign n568 = ~n566 & ~n567;
  assign n569 = n565 & ~n568;
  assign n570 = ~n565 & n568;
  assign \f[23]  = ~n569 & ~n570;
  assign n572 = ~n565 & ~n566;
  assign n573 = ~n567 & ~n572;
  assign n574 = ~\a[24]  & ~\b[24] ;
  assign n575 = \a[24]  & \b[24] ;
  assign n576 = ~n574 & ~n575;
  assign n577 = n573 & ~n576;
  assign n578 = ~n573 & n576;
  assign \f[24]  = ~n577 & ~n578;
  assign n580 = ~n573 & ~n574;
  assign n581 = ~n575 & ~n580;
  assign n582 = ~\a[25]  & ~\b[25] ;
  assign n583 = \a[25]  & \b[25] ;
  assign n584 = ~n582 & ~n583;
  assign n585 = n581 & ~n584;
  assign n586 = ~n581 & n584;
  assign \f[25]  = ~n585 & ~n586;
  assign n588 = ~n581 & ~n582;
  assign n589 = ~n583 & ~n588;
  assign n590 = ~\a[26]  & ~\b[26] ;
  assign n591 = \a[26]  & \b[26] ;
  assign n592 = ~n590 & ~n591;
  assign n593 = n589 & ~n592;
  assign n594 = ~n589 & n592;
  assign \f[26]  = ~n593 & ~n594;
  assign n596 = ~n589 & ~n590;
  assign n597 = ~n591 & ~n596;
  assign n598 = ~\a[27]  & ~\b[27] ;
  assign n599 = \a[27]  & \b[27] ;
  assign n600 = ~n598 & ~n599;
  assign n601 = n597 & ~n600;
  assign n602 = ~n597 & n600;
  assign \f[27]  = ~n601 & ~n602;
  assign n604 = ~n597 & ~n598;
  assign n605 = ~n599 & ~n604;
  assign n606 = ~\a[28]  & ~\b[28] ;
  assign n607 = \a[28]  & \b[28] ;
  assign n608 = ~n606 & ~n607;
  assign n609 = n605 & ~n608;
  assign n610 = ~n605 & n608;
  assign \f[28]  = ~n609 & ~n610;
  assign n612 = ~n605 & ~n606;
  assign n613 = ~n607 & ~n612;
  assign n614 = ~\a[29]  & ~\b[29] ;
  assign n615 = \a[29]  & \b[29] ;
  assign n616 = ~n614 & ~n615;
  assign n617 = n613 & ~n616;
  assign n618 = ~n613 & n616;
  assign \f[29]  = ~n617 & ~n618;
  assign n620 = ~n613 & ~n614;
  assign n621 = ~n615 & ~n620;
  assign n622 = ~\a[30]  & ~\b[30] ;
  assign n623 = \a[30]  & \b[30] ;
  assign n624 = ~n622 & ~n623;
  assign n625 = n621 & ~n624;
  assign n626 = ~n621 & n624;
  assign \f[30]  = ~n625 & ~n626;
  assign n628 = ~n621 & ~n622;
  assign n629 = ~n623 & ~n628;
  assign n630 = ~\a[31]  & ~\b[31] ;
  assign n631 = \a[31]  & \b[31] ;
  assign n632 = ~n630 & ~n631;
  assign n633 = n629 & ~n632;
  assign n634 = ~n629 & n632;
  assign \f[31]  = ~n633 & ~n634;
  assign n636 = ~n629 & ~n630;
  assign n637 = ~n631 & ~n636;
  assign n638 = ~\a[32]  & ~\b[32] ;
  assign n639 = \a[32]  & \b[32] ;
  assign n640 = ~n638 & ~n639;
  assign n641 = n637 & ~n640;
  assign n642 = ~n637 & n640;
  assign \f[32]  = ~n641 & ~n642;
  assign n644 = ~n637 & ~n638;
  assign n645 = ~n639 & ~n644;
  assign n646 = ~\a[33]  & ~\b[33] ;
  assign n647 = \a[33]  & \b[33] ;
  assign n648 = ~n646 & ~n647;
  assign n649 = n645 & ~n648;
  assign n650 = ~n645 & n648;
  assign \f[33]  = ~n649 & ~n650;
  assign n652 = ~n645 & ~n646;
  assign n653 = ~n647 & ~n652;
  assign n654 = ~\a[34]  & ~\b[34] ;
  assign n655 = \a[34]  & \b[34] ;
  assign n656 = ~n654 & ~n655;
  assign n657 = n653 & ~n656;
  assign n658 = ~n653 & n656;
  assign \f[34]  = ~n657 & ~n658;
  assign n660 = ~n653 & ~n654;
  assign n661 = ~n655 & ~n660;
  assign n662 = ~\a[35]  & ~\b[35] ;
  assign n663 = \a[35]  & \b[35] ;
  assign n664 = ~n662 & ~n663;
  assign n665 = n661 & ~n664;
  assign n666 = ~n661 & n664;
  assign \f[35]  = ~n665 & ~n666;
  assign n668 = ~n661 & ~n662;
  assign n669 = ~n663 & ~n668;
  assign n670 = ~\a[36]  & ~\b[36] ;
  assign n671 = \a[36]  & \b[36] ;
  assign n672 = ~n670 & ~n671;
  assign n673 = n669 & ~n672;
  assign n674 = ~n669 & n672;
  assign \f[36]  = ~n673 & ~n674;
  assign n676 = ~n669 & ~n670;
  assign n677 = ~n671 & ~n676;
  assign n678 = ~\a[37]  & ~\b[37] ;
  assign n679 = \a[37]  & \b[37] ;
  assign n680 = ~n678 & ~n679;
  assign n681 = n677 & ~n680;
  assign n682 = ~n677 & n680;
  assign \f[37]  = ~n681 & ~n682;
  assign n684 = ~n677 & ~n678;
  assign n685 = ~n679 & ~n684;
  assign n686 = ~\a[38]  & ~\b[38] ;
  assign n687 = \a[38]  & \b[38] ;
  assign n688 = ~n686 & ~n687;
  assign n689 = n685 & ~n688;
  assign n690 = ~n685 & n688;
  assign \f[38]  = ~n689 & ~n690;
  assign n692 = ~n685 & ~n686;
  assign n693 = ~n687 & ~n692;
  assign n694 = ~\a[39]  & ~\b[39] ;
  assign n695 = \a[39]  & \b[39] ;
  assign n696 = ~n694 & ~n695;
  assign n697 = n693 & ~n696;
  assign n698 = ~n693 & n696;
  assign \f[39]  = ~n697 & ~n698;
  assign n700 = ~n693 & ~n694;
  assign n701 = ~n695 & ~n700;
  assign n702 = ~\a[40]  & ~\b[40] ;
  assign n703 = \a[40]  & \b[40] ;
  assign n704 = ~n702 & ~n703;
  assign n705 = n701 & ~n704;
  assign n706 = ~n701 & n704;
  assign \f[40]  = ~n705 & ~n706;
  assign n708 = ~n701 & ~n702;
  assign n709 = ~n703 & ~n708;
  assign n710 = ~\a[41]  & ~\b[41] ;
  assign n711 = \a[41]  & \b[41] ;
  assign n712 = ~n710 & ~n711;
  assign n713 = n709 & ~n712;
  assign n714 = ~n709 & n712;
  assign \f[41]  = ~n713 & ~n714;
  assign n716 = ~n709 & ~n710;
  assign n717 = ~n711 & ~n716;
  assign n718 = ~\a[42]  & ~\b[42] ;
  assign n719 = \a[42]  & \b[42] ;
  assign n720 = ~n718 & ~n719;
  assign n721 = n717 & ~n720;
  assign n722 = ~n717 & n720;
  assign \f[42]  = ~n721 & ~n722;
  assign n724 = ~n717 & ~n718;
  assign n725 = ~n719 & ~n724;
  assign n726 = ~\a[43]  & ~\b[43] ;
  assign n727 = \a[43]  & \b[43] ;
  assign n728 = ~n726 & ~n727;
  assign n729 = n725 & ~n728;
  assign n730 = ~n725 & n728;
  assign \f[43]  = ~n729 & ~n730;
  assign n732 = ~n725 & ~n726;
  assign n733 = ~n727 & ~n732;
  assign n734 = ~\a[44]  & ~\b[44] ;
  assign n735 = \a[44]  & \b[44] ;
  assign n736 = ~n734 & ~n735;
  assign n737 = n733 & ~n736;
  assign n738 = ~n733 & n736;
  assign \f[44]  = ~n737 & ~n738;
  assign n740 = ~n733 & ~n734;
  assign n741 = ~n735 & ~n740;
  assign n742 = ~\a[45]  & ~\b[45] ;
  assign n743 = \a[45]  & \b[45] ;
  assign n744 = ~n742 & ~n743;
  assign n745 = n741 & ~n744;
  assign n746 = ~n741 & n744;
  assign \f[45]  = ~n745 & ~n746;
  assign n748 = ~n741 & ~n742;
  assign n749 = ~n743 & ~n748;
  assign n750 = ~\a[46]  & ~\b[46] ;
  assign n751 = \a[46]  & \b[46] ;
  assign n752 = ~n750 & ~n751;
  assign n753 = n749 & ~n752;
  assign n754 = ~n749 & n752;
  assign \f[46]  = ~n753 & ~n754;
  assign n756 = ~n749 & ~n750;
  assign n757 = ~n751 & ~n756;
  assign n758 = ~\a[47]  & ~\b[47] ;
  assign n759 = \a[47]  & \b[47] ;
  assign n760 = ~n758 & ~n759;
  assign n761 = n757 & ~n760;
  assign n762 = ~n757 & n760;
  assign \f[47]  = ~n761 & ~n762;
  assign n764 = ~n757 & ~n758;
  assign n765 = ~n759 & ~n764;
  assign n766 = ~\a[48]  & ~\b[48] ;
  assign n767 = \a[48]  & \b[48] ;
  assign n768 = ~n766 & ~n767;
  assign n769 = n765 & ~n768;
  assign n770 = ~n765 & n768;
  assign \f[48]  = ~n769 & ~n770;
  assign n772 = ~n765 & ~n766;
  assign n773 = ~n767 & ~n772;
  assign n774 = ~\a[49]  & ~\b[49] ;
  assign n775 = \a[49]  & \b[49] ;
  assign n776 = ~n774 & ~n775;
  assign n777 = n773 & ~n776;
  assign n778 = ~n773 & n776;
  assign \f[49]  = ~n777 & ~n778;
  assign n780 = ~n773 & ~n774;
  assign n781 = ~n775 & ~n780;
  assign n782 = ~\a[50]  & ~\b[50] ;
  assign n783 = \a[50]  & \b[50] ;
  assign n784 = ~n782 & ~n783;
  assign n785 = n781 & ~n784;
  assign n786 = ~n781 & n784;
  assign \f[50]  = ~n785 & ~n786;
  assign n788 = ~n781 & ~n782;
  assign n789 = ~n783 & ~n788;
  assign n790 = ~\a[51]  & ~\b[51] ;
  assign n791 = \a[51]  & \b[51] ;
  assign n792 = ~n790 & ~n791;
  assign n793 = n789 & ~n792;
  assign n794 = ~n789 & n792;
  assign \f[51]  = ~n793 & ~n794;
  assign n796 = ~n789 & ~n790;
  assign n797 = ~n791 & ~n796;
  assign n798 = ~\a[52]  & ~\b[52] ;
  assign n799 = \a[52]  & \b[52] ;
  assign n800 = ~n798 & ~n799;
  assign n801 = n797 & ~n800;
  assign n802 = ~n797 & n800;
  assign \f[52]  = ~n801 & ~n802;
  assign n804 = ~n797 & ~n798;
  assign n805 = ~n799 & ~n804;
  assign n806 = ~\a[53]  & ~\b[53] ;
  assign n807 = \a[53]  & \b[53] ;
  assign n808 = ~n806 & ~n807;
  assign n809 = n805 & ~n808;
  assign n810 = ~n805 & n808;
  assign \f[53]  = ~n809 & ~n810;
  assign n812 = ~n805 & ~n806;
  assign n813 = ~n807 & ~n812;
  assign n814 = ~\a[54]  & ~\b[54] ;
  assign n815 = \a[54]  & \b[54] ;
  assign n816 = ~n814 & ~n815;
  assign n817 = n813 & ~n816;
  assign n818 = ~n813 & n816;
  assign \f[54]  = ~n817 & ~n818;
  assign n820 = ~n813 & ~n814;
  assign n821 = ~n815 & ~n820;
  assign n822 = ~\a[55]  & ~\b[55] ;
  assign n823 = \a[55]  & \b[55] ;
  assign n824 = ~n822 & ~n823;
  assign n825 = n821 & ~n824;
  assign n826 = ~n821 & n824;
  assign \f[55]  = ~n825 & ~n826;
  assign n828 = ~n821 & ~n822;
  assign n829 = ~n823 & ~n828;
  assign n830 = ~\a[56]  & ~\b[56] ;
  assign n831 = \a[56]  & \b[56] ;
  assign n832 = ~n830 & ~n831;
  assign n833 = n829 & ~n832;
  assign n834 = ~n829 & n832;
  assign \f[56]  = ~n833 & ~n834;
  assign n836 = ~n829 & ~n830;
  assign n837 = ~n831 & ~n836;
  assign n838 = ~\a[57]  & ~\b[57] ;
  assign n839 = \a[57]  & \b[57] ;
  assign n840 = ~n838 & ~n839;
  assign n841 = n837 & ~n840;
  assign n842 = ~n837 & n840;
  assign \f[57]  = ~n841 & ~n842;
  assign n844 = ~n837 & ~n838;
  assign n845 = ~n839 & ~n844;
  assign n846 = ~\a[58]  & ~\b[58] ;
  assign n847 = \a[58]  & \b[58] ;
  assign n848 = ~n846 & ~n847;
  assign n849 = n845 & ~n848;
  assign n850 = ~n845 & n848;
  assign \f[58]  = ~n849 & ~n850;
  assign n852 = ~n845 & ~n846;
  assign n853 = ~n847 & ~n852;
  assign n854 = ~\a[59]  & ~\b[59] ;
  assign n855 = \a[59]  & \b[59] ;
  assign n856 = ~n854 & ~n855;
  assign n857 = n853 & ~n856;
  assign n858 = ~n853 & n856;
  assign \f[59]  = ~n857 & ~n858;
  assign n860 = ~n853 & ~n854;
  assign n861 = ~n855 & ~n860;
  assign n862 = ~\a[60]  & ~\b[60] ;
  assign n863 = \a[60]  & \b[60] ;
  assign n864 = ~n862 & ~n863;
  assign n865 = n861 & ~n864;
  assign n866 = ~n861 & n864;
  assign \f[60]  = ~n865 & ~n866;
  assign n868 = ~n861 & ~n862;
  assign n869 = ~n863 & ~n868;
  assign n870 = ~\a[61]  & ~\b[61] ;
  assign n871 = \a[61]  & \b[61] ;
  assign n872 = ~n870 & ~n871;
  assign n873 = n869 & ~n872;
  assign n874 = ~n869 & n872;
  assign \f[61]  = ~n873 & ~n874;
  assign n876 = ~n869 & ~n870;
  assign n877 = ~n871 & ~n876;
  assign n878 = ~\a[62]  & ~\b[62] ;
  assign n879 = \a[62]  & \b[62] ;
  assign n880 = ~n878 & ~n879;
  assign n881 = n877 & ~n880;
  assign n882 = ~n877 & n880;
  assign \f[62]  = ~n881 & ~n882;
  assign n884 = ~n877 & ~n878;
  assign n885 = ~n879 & ~n884;
  assign n886 = ~\a[63]  & ~\b[63] ;
  assign n887 = \a[63]  & \b[63] ;
  assign n888 = ~n886 & ~n887;
  assign n889 = n885 & ~n888;
  assign n890 = ~n885 & n888;
  assign \f[63]  = ~n889 & ~n890;
  assign n892 = ~n885 & ~n886;
  assign n893 = ~n887 & ~n892;
  assign n894 = ~\a[64]  & ~\b[64] ;
  assign n895 = \a[64]  & \b[64] ;
  assign n896 = ~n894 & ~n895;
  assign n897 = n893 & ~n896;
  assign n898 = ~n893 & n896;
  assign \f[64]  = ~n897 & ~n898;
  assign n900 = ~n893 & ~n894;
  assign n901 = ~n895 & ~n900;
  assign n902 = ~\a[65]  & ~\b[65] ;
  assign n903 = \a[65]  & \b[65] ;
  assign n904 = ~n902 & ~n903;
  assign n905 = n901 & ~n904;
  assign n906 = ~n901 & n904;
  assign \f[65]  = ~n905 & ~n906;
  assign n908 = ~n901 & ~n902;
  assign n909 = ~n903 & ~n908;
  assign n910 = ~\a[66]  & ~\b[66] ;
  assign n911 = \a[66]  & \b[66] ;
  assign n912 = ~n910 & ~n911;
  assign n913 = n909 & ~n912;
  assign n914 = ~n909 & n912;
  assign \f[66]  = ~n913 & ~n914;
  assign n916 = ~n909 & ~n910;
  assign n917 = ~n911 & ~n916;
  assign n918 = ~\a[67]  & ~\b[67] ;
  assign n919 = \a[67]  & \b[67] ;
  assign n920 = ~n918 & ~n919;
  assign n921 = n917 & ~n920;
  assign n922 = ~n917 & n920;
  assign \f[67]  = ~n921 & ~n922;
  assign n924 = ~n917 & ~n918;
  assign n925 = ~n919 & ~n924;
  assign n926 = ~\a[68]  & ~\b[68] ;
  assign n927 = \a[68]  & \b[68] ;
  assign n928 = ~n926 & ~n927;
  assign n929 = n925 & ~n928;
  assign n930 = ~n925 & n928;
  assign \f[68]  = ~n929 & ~n930;
  assign n932 = ~n925 & ~n926;
  assign n933 = ~n927 & ~n932;
  assign n934 = ~\a[69]  & ~\b[69] ;
  assign n935 = \a[69]  & \b[69] ;
  assign n936 = ~n934 & ~n935;
  assign n937 = n933 & ~n936;
  assign n938 = ~n933 & n936;
  assign \f[69]  = ~n937 & ~n938;
  assign n940 = ~n933 & ~n934;
  assign n941 = ~n935 & ~n940;
  assign n942 = ~\a[70]  & ~\b[70] ;
  assign n943 = \a[70]  & \b[70] ;
  assign n944 = ~n942 & ~n943;
  assign n945 = n941 & ~n944;
  assign n946 = ~n941 & n944;
  assign \f[70]  = ~n945 & ~n946;
  assign n948 = ~n941 & ~n942;
  assign n949 = ~n943 & ~n948;
  assign n950 = ~\a[71]  & ~\b[71] ;
  assign n951 = \a[71]  & \b[71] ;
  assign n952 = ~n950 & ~n951;
  assign n953 = n949 & ~n952;
  assign n954 = ~n949 & n952;
  assign \f[71]  = ~n953 & ~n954;
  assign n956 = ~n949 & ~n950;
  assign n957 = ~n951 & ~n956;
  assign n958 = ~\a[72]  & ~\b[72] ;
  assign n959 = \a[72]  & \b[72] ;
  assign n960 = ~n958 & ~n959;
  assign n961 = n957 & ~n960;
  assign n962 = ~n957 & n960;
  assign \f[72]  = ~n961 & ~n962;
  assign n964 = ~n957 & ~n958;
  assign n965 = ~n959 & ~n964;
  assign n966 = ~\a[73]  & ~\b[73] ;
  assign n967 = \a[73]  & \b[73] ;
  assign n968 = ~n966 & ~n967;
  assign n969 = n965 & ~n968;
  assign n970 = ~n965 & n968;
  assign \f[73]  = ~n969 & ~n970;
  assign n972 = ~n965 & ~n966;
  assign n973 = ~n967 & ~n972;
  assign n974 = ~\a[74]  & ~\b[74] ;
  assign n975 = \a[74]  & \b[74] ;
  assign n976 = ~n974 & ~n975;
  assign n977 = n973 & ~n976;
  assign n978 = ~n973 & n976;
  assign \f[74]  = ~n977 & ~n978;
  assign n980 = ~n973 & ~n974;
  assign n981 = ~n975 & ~n980;
  assign n982 = ~\a[75]  & ~\b[75] ;
  assign n983 = \a[75]  & \b[75] ;
  assign n984 = ~n982 & ~n983;
  assign n985 = n981 & ~n984;
  assign n986 = ~n981 & n984;
  assign \f[75]  = ~n985 & ~n986;
  assign n988 = ~n981 & ~n982;
  assign n989 = ~n983 & ~n988;
  assign n990 = ~\a[76]  & ~\b[76] ;
  assign n991 = \a[76]  & \b[76] ;
  assign n992 = ~n990 & ~n991;
  assign n993 = n989 & ~n992;
  assign n994 = ~n989 & n992;
  assign \f[76]  = ~n993 & ~n994;
  assign n996 = ~n989 & ~n990;
  assign n997 = ~n991 & ~n996;
  assign n998 = ~\a[77]  & ~\b[77] ;
  assign n999 = \a[77]  & \b[77] ;
  assign n1000 = ~n998 & ~n999;
  assign n1001 = n997 & ~n1000;
  assign n1002 = ~n997 & n1000;
  assign \f[77]  = ~n1001 & ~n1002;
  assign n1004 = ~n997 & ~n998;
  assign n1005 = ~n999 & ~n1004;
  assign n1006 = ~\a[78]  & ~\b[78] ;
  assign n1007 = \a[78]  & \b[78] ;
  assign n1008 = ~n1006 & ~n1007;
  assign n1009 = n1005 & ~n1008;
  assign n1010 = ~n1005 & n1008;
  assign \f[78]  = ~n1009 & ~n1010;
  assign n1012 = ~n1005 & ~n1006;
  assign n1013 = ~n1007 & ~n1012;
  assign n1014 = ~\a[79]  & ~\b[79] ;
  assign n1015 = \a[79]  & \b[79] ;
  assign n1016 = ~n1014 & ~n1015;
  assign n1017 = n1013 & ~n1016;
  assign n1018 = ~n1013 & n1016;
  assign \f[79]  = ~n1017 & ~n1018;
  assign n1020 = ~n1013 & ~n1014;
  assign n1021 = ~n1015 & ~n1020;
  assign n1022 = ~\a[80]  & ~\b[80] ;
  assign n1023 = \a[80]  & \b[80] ;
  assign n1024 = ~n1022 & ~n1023;
  assign n1025 = n1021 & ~n1024;
  assign n1026 = ~n1021 & n1024;
  assign \f[80]  = ~n1025 & ~n1026;
  assign n1028 = ~n1021 & ~n1022;
  assign n1029 = ~n1023 & ~n1028;
  assign n1030 = ~\a[81]  & ~\b[81] ;
  assign n1031 = \a[81]  & \b[81] ;
  assign n1032 = ~n1030 & ~n1031;
  assign n1033 = n1029 & ~n1032;
  assign n1034 = ~n1029 & n1032;
  assign \f[81]  = ~n1033 & ~n1034;
  assign n1036 = ~n1029 & ~n1030;
  assign n1037 = ~n1031 & ~n1036;
  assign n1038 = ~\a[82]  & ~\b[82] ;
  assign n1039 = \a[82]  & \b[82] ;
  assign n1040 = ~n1038 & ~n1039;
  assign n1041 = n1037 & ~n1040;
  assign n1042 = ~n1037 & n1040;
  assign \f[82]  = ~n1041 & ~n1042;
  assign n1044 = ~n1037 & ~n1038;
  assign n1045 = ~n1039 & ~n1044;
  assign n1046 = ~\a[83]  & ~\b[83] ;
  assign n1047 = \a[83]  & \b[83] ;
  assign n1048 = ~n1046 & ~n1047;
  assign n1049 = n1045 & ~n1048;
  assign n1050 = ~n1045 & n1048;
  assign \f[83]  = ~n1049 & ~n1050;
  assign n1052 = ~n1045 & ~n1046;
  assign n1053 = ~n1047 & ~n1052;
  assign n1054 = ~\a[84]  & ~\b[84] ;
  assign n1055 = \a[84]  & \b[84] ;
  assign n1056 = ~n1054 & ~n1055;
  assign n1057 = n1053 & ~n1056;
  assign n1058 = ~n1053 & n1056;
  assign \f[84]  = ~n1057 & ~n1058;
  assign n1060 = ~n1053 & ~n1054;
  assign n1061 = ~n1055 & ~n1060;
  assign n1062 = ~\a[85]  & ~\b[85] ;
  assign n1063 = \a[85]  & \b[85] ;
  assign n1064 = ~n1062 & ~n1063;
  assign n1065 = n1061 & ~n1064;
  assign n1066 = ~n1061 & n1064;
  assign \f[85]  = ~n1065 & ~n1066;
  assign n1068 = ~n1061 & ~n1062;
  assign n1069 = ~n1063 & ~n1068;
  assign n1070 = ~\a[86]  & ~\b[86] ;
  assign n1071 = \a[86]  & \b[86] ;
  assign n1072 = ~n1070 & ~n1071;
  assign n1073 = n1069 & ~n1072;
  assign n1074 = ~n1069 & n1072;
  assign \f[86]  = ~n1073 & ~n1074;
  assign n1076 = ~n1069 & ~n1070;
  assign n1077 = ~n1071 & ~n1076;
  assign n1078 = ~\a[87]  & ~\b[87] ;
  assign n1079 = \a[87]  & \b[87] ;
  assign n1080 = ~n1078 & ~n1079;
  assign n1081 = n1077 & ~n1080;
  assign n1082 = ~n1077 & n1080;
  assign \f[87]  = ~n1081 & ~n1082;
  assign n1084 = ~n1077 & ~n1078;
  assign n1085 = ~n1079 & ~n1084;
  assign n1086 = ~\a[88]  & ~\b[88] ;
  assign n1087 = \a[88]  & \b[88] ;
  assign n1088 = ~n1086 & ~n1087;
  assign n1089 = n1085 & ~n1088;
  assign n1090 = ~n1085 & n1088;
  assign \f[88]  = ~n1089 & ~n1090;
  assign n1092 = ~n1085 & ~n1086;
  assign n1093 = ~n1087 & ~n1092;
  assign n1094 = ~\a[89]  & ~\b[89] ;
  assign n1095 = \a[89]  & \b[89] ;
  assign n1096 = ~n1094 & ~n1095;
  assign n1097 = n1093 & ~n1096;
  assign n1098 = ~n1093 & n1096;
  assign \f[89]  = ~n1097 & ~n1098;
  assign n1100 = ~n1093 & ~n1094;
  assign n1101 = ~n1095 & ~n1100;
  assign n1102 = ~\a[90]  & ~\b[90] ;
  assign n1103 = \a[90]  & \b[90] ;
  assign n1104 = ~n1102 & ~n1103;
  assign n1105 = n1101 & ~n1104;
  assign n1106 = ~n1101 & n1104;
  assign \f[90]  = ~n1105 & ~n1106;
  assign n1108 = ~n1101 & ~n1102;
  assign n1109 = ~n1103 & ~n1108;
  assign n1110 = ~\a[91]  & ~\b[91] ;
  assign n1111 = \a[91]  & \b[91] ;
  assign n1112 = ~n1110 & ~n1111;
  assign n1113 = n1109 & ~n1112;
  assign n1114 = ~n1109 & n1112;
  assign \f[91]  = ~n1113 & ~n1114;
  assign n1116 = ~n1109 & ~n1110;
  assign n1117 = ~n1111 & ~n1116;
  assign n1118 = ~\a[92]  & ~\b[92] ;
  assign n1119 = \a[92]  & \b[92] ;
  assign n1120 = ~n1118 & ~n1119;
  assign n1121 = n1117 & ~n1120;
  assign n1122 = ~n1117 & n1120;
  assign \f[92]  = ~n1121 & ~n1122;
  assign n1124 = ~n1117 & ~n1118;
  assign n1125 = ~n1119 & ~n1124;
  assign n1126 = ~\a[93]  & ~\b[93] ;
  assign n1127 = \a[93]  & \b[93] ;
  assign n1128 = ~n1126 & ~n1127;
  assign n1129 = n1125 & ~n1128;
  assign n1130 = ~n1125 & n1128;
  assign \f[93]  = ~n1129 & ~n1130;
  assign n1132 = ~n1125 & ~n1126;
  assign n1133 = ~n1127 & ~n1132;
  assign n1134 = ~\a[94]  & ~\b[94] ;
  assign n1135 = \a[94]  & \b[94] ;
  assign n1136 = ~n1134 & ~n1135;
  assign n1137 = n1133 & ~n1136;
  assign n1138 = ~n1133 & n1136;
  assign \f[94]  = ~n1137 & ~n1138;
  assign n1140 = ~n1133 & ~n1134;
  assign n1141 = ~n1135 & ~n1140;
  assign n1142 = ~\a[95]  & ~\b[95] ;
  assign n1143 = \a[95]  & \b[95] ;
  assign n1144 = ~n1142 & ~n1143;
  assign n1145 = n1141 & ~n1144;
  assign n1146 = ~n1141 & n1144;
  assign \f[95]  = ~n1145 & ~n1146;
  assign n1148 = ~n1141 & ~n1142;
  assign n1149 = ~n1143 & ~n1148;
  assign n1150 = ~\a[96]  & ~\b[96] ;
  assign n1151 = \a[96]  & \b[96] ;
  assign n1152 = ~n1150 & ~n1151;
  assign n1153 = n1149 & ~n1152;
  assign n1154 = ~n1149 & n1152;
  assign \f[96]  = ~n1153 & ~n1154;
  assign n1156 = ~n1149 & ~n1150;
  assign n1157 = ~n1151 & ~n1156;
  assign n1158 = ~\a[97]  & ~\b[97] ;
  assign n1159 = \a[97]  & \b[97] ;
  assign n1160 = ~n1158 & ~n1159;
  assign n1161 = n1157 & ~n1160;
  assign n1162 = ~n1157 & n1160;
  assign \f[97]  = ~n1161 & ~n1162;
  assign n1164 = ~n1157 & ~n1158;
  assign n1165 = ~n1159 & ~n1164;
  assign n1166 = ~\a[98]  & ~\b[98] ;
  assign n1167 = \a[98]  & \b[98] ;
  assign n1168 = ~n1166 & ~n1167;
  assign n1169 = n1165 & ~n1168;
  assign n1170 = ~n1165 & n1168;
  assign \f[98]  = ~n1169 & ~n1170;
  assign n1172 = ~n1165 & ~n1166;
  assign n1173 = ~n1167 & ~n1172;
  assign n1174 = ~\a[99]  & ~\b[99] ;
  assign n1175 = \a[99]  & \b[99] ;
  assign n1176 = ~n1174 & ~n1175;
  assign n1177 = n1173 & ~n1176;
  assign n1178 = ~n1173 & n1176;
  assign \f[99]  = ~n1177 & ~n1178;
  assign n1180 = ~n1173 & ~n1174;
  assign n1181 = ~n1175 & ~n1180;
  assign n1182 = ~\a[100]  & ~\b[100] ;
  assign n1183 = \a[100]  & \b[100] ;
  assign n1184 = ~n1182 & ~n1183;
  assign n1185 = n1181 & ~n1184;
  assign n1186 = ~n1181 & n1184;
  assign \f[100]  = ~n1185 & ~n1186;
  assign n1188 = ~n1181 & ~n1182;
  assign n1189 = ~n1183 & ~n1188;
  assign n1190 = ~\a[101]  & ~\b[101] ;
  assign n1191 = \a[101]  & \b[101] ;
  assign n1192 = ~n1190 & ~n1191;
  assign n1193 = n1189 & ~n1192;
  assign n1194 = ~n1189 & n1192;
  assign \f[101]  = ~n1193 & ~n1194;
  assign n1196 = ~n1189 & ~n1190;
  assign n1197 = ~n1191 & ~n1196;
  assign n1198 = ~\a[102]  & ~\b[102] ;
  assign n1199 = \a[102]  & \b[102] ;
  assign n1200 = ~n1198 & ~n1199;
  assign n1201 = n1197 & ~n1200;
  assign n1202 = ~n1197 & n1200;
  assign \f[102]  = ~n1201 & ~n1202;
  assign n1204 = ~n1197 & ~n1198;
  assign n1205 = ~n1199 & ~n1204;
  assign n1206 = ~\a[103]  & ~\b[103] ;
  assign n1207 = \a[103]  & \b[103] ;
  assign n1208 = ~n1206 & ~n1207;
  assign n1209 = n1205 & ~n1208;
  assign n1210 = ~n1205 & n1208;
  assign \f[103]  = ~n1209 & ~n1210;
  assign n1212 = ~n1205 & ~n1206;
  assign n1213 = ~n1207 & ~n1212;
  assign n1214 = ~\a[104]  & ~\b[104] ;
  assign n1215 = \a[104]  & \b[104] ;
  assign n1216 = ~n1214 & ~n1215;
  assign n1217 = n1213 & ~n1216;
  assign n1218 = ~n1213 & n1216;
  assign \f[104]  = ~n1217 & ~n1218;
  assign n1220 = ~n1213 & ~n1214;
  assign n1221 = ~n1215 & ~n1220;
  assign n1222 = ~\a[105]  & ~\b[105] ;
  assign n1223 = \a[105]  & \b[105] ;
  assign n1224 = ~n1222 & ~n1223;
  assign n1225 = n1221 & ~n1224;
  assign n1226 = ~n1221 & n1224;
  assign \f[105]  = ~n1225 & ~n1226;
  assign n1228 = ~n1221 & ~n1222;
  assign n1229 = ~n1223 & ~n1228;
  assign n1230 = ~\a[106]  & ~\b[106] ;
  assign n1231 = \a[106]  & \b[106] ;
  assign n1232 = ~n1230 & ~n1231;
  assign n1233 = n1229 & ~n1232;
  assign n1234 = ~n1229 & n1232;
  assign \f[106]  = ~n1233 & ~n1234;
  assign n1236 = ~n1229 & ~n1230;
  assign n1237 = ~n1231 & ~n1236;
  assign n1238 = ~\a[107]  & ~\b[107] ;
  assign n1239 = \a[107]  & \b[107] ;
  assign n1240 = ~n1238 & ~n1239;
  assign n1241 = n1237 & ~n1240;
  assign n1242 = ~n1237 & n1240;
  assign \f[107]  = ~n1241 & ~n1242;
  assign n1244 = ~n1237 & ~n1238;
  assign n1245 = ~n1239 & ~n1244;
  assign n1246 = ~\a[108]  & ~\b[108] ;
  assign n1247 = \a[108]  & \b[108] ;
  assign n1248 = ~n1246 & ~n1247;
  assign n1249 = n1245 & ~n1248;
  assign n1250 = ~n1245 & n1248;
  assign \f[108]  = ~n1249 & ~n1250;
  assign n1252 = ~n1245 & ~n1246;
  assign n1253 = ~n1247 & ~n1252;
  assign n1254 = ~\a[109]  & ~\b[109] ;
  assign n1255 = \a[109]  & \b[109] ;
  assign n1256 = ~n1254 & ~n1255;
  assign n1257 = n1253 & ~n1256;
  assign n1258 = ~n1253 & n1256;
  assign \f[109]  = ~n1257 & ~n1258;
  assign n1260 = ~n1253 & ~n1254;
  assign n1261 = ~n1255 & ~n1260;
  assign n1262 = ~\a[110]  & ~\b[110] ;
  assign n1263 = \a[110]  & \b[110] ;
  assign n1264 = ~n1262 & ~n1263;
  assign n1265 = n1261 & ~n1264;
  assign n1266 = ~n1261 & n1264;
  assign \f[110]  = ~n1265 & ~n1266;
  assign n1268 = ~n1261 & ~n1262;
  assign n1269 = ~n1263 & ~n1268;
  assign n1270 = ~\a[111]  & ~\b[111] ;
  assign n1271 = \a[111]  & \b[111] ;
  assign n1272 = ~n1270 & ~n1271;
  assign n1273 = n1269 & ~n1272;
  assign n1274 = ~n1269 & n1272;
  assign \f[111]  = ~n1273 & ~n1274;
  assign n1276 = ~n1269 & ~n1270;
  assign n1277 = ~n1271 & ~n1276;
  assign n1278 = ~\a[112]  & ~\b[112] ;
  assign n1279 = \a[112]  & \b[112] ;
  assign n1280 = ~n1278 & ~n1279;
  assign n1281 = n1277 & ~n1280;
  assign n1282 = ~n1277 & n1280;
  assign \f[112]  = ~n1281 & ~n1282;
  assign n1284 = ~n1277 & ~n1278;
  assign n1285 = ~n1279 & ~n1284;
  assign n1286 = ~\a[113]  & ~\b[113] ;
  assign n1287 = \a[113]  & \b[113] ;
  assign n1288 = ~n1286 & ~n1287;
  assign n1289 = n1285 & ~n1288;
  assign n1290 = ~n1285 & n1288;
  assign \f[113]  = ~n1289 & ~n1290;
  assign n1292 = ~n1285 & ~n1286;
  assign n1293 = ~n1287 & ~n1292;
  assign n1294 = ~\a[114]  & ~\b[114] ;
  assign n1295 = \a[114]  & \b[114] ;
  assign n1296 = ~n1294 & ~n1295;
  assign n1297 = n1293 & ~n1296;
  assign n1298 = ~n1293 & n1296;
  assign \f[114]  = ~n1297 & ~n1298;
  assign n1300 = ~n1293 & ~n1294;
  assign n1301 = ~n1295 & ~n1300;
  assign n1302 = ~\a[115]  & ~\b[115] ;
  assign n1303 = \a[115]  & \b[115] ;
  assign n1304 = ~n1302 & ~n1303;
  assign n1305 = n1301 & ~n1304;
  assign n1306 = ~n1301 & n1304;
  assign \f[115]  = ~n1305 & ~n1306;
  assign n1308 = ~n1301 & ~n1302;
  assign n1309 = ~n1303 & ~n1308;
  assign n1310 = ~\a[116]  & ~\b[116] ;
  assign n1311 = \a[116]  & \b[116] ;
  assign n1312 = ~n1310 & ~n1311;
  assign n1313 = n1309 & ~n1312;
  assign n1314 = ~n1309 & n1312;
  assign \f[116]  = ~n1313 & ~n1314;
  assign n1316 = ~n1309 & ~n1310;
  assign n1317 = ~n1311 & ~n1316;
  assign n1318 = ~\a[117]  & ~\b[117] ;
  assign n1319 = \a[117]  & \b[117] ;
  assign n1320 = ~n1318 & ~n1319;
  assign n1321 = n1317 & ~n1320;
  assign n1322 = ~n1317 & n1320;
  assign \f[117]  = ~n1321 & ~n1322;
  assign n1324 = ~n1317 & ~n1318;
  assign n1325 = ~n1319 & ~n1324;
  assign n1326 = ~\a[118]  & ~\b[118] ;
  assign n1327 = \a[118]  & \b[118] ;
  assign n1328 = ~n1326 & ~n1327;
  assign n1329 = n1325 & ~n1328;
  assign n1330 = ~n1325 & n1328;
  assign \f[118]  = ~n1329 & ~n1330;
  assign n1332 = ~n1325 & ~n1326;
  assign n1333 = ~n1327 & ~n1332;
  assign n1334 = ~\a[119]  & ~\b[119] ;
  assign n1335 = \a[119]  & \b[119] ;
  assign n1336 = ~n1334 & ~n1335;
  assign n1337 = n1333 & ~n1336;
  assign n1338 = ~n1333 & n1336;
  assign \f[119]  = ~n1337 & ~n1338;
  assign n1340 = ~n1333 & ~n1334;
  assign n1341 = ~n1335 & ~n1340;
  assign n1342 = ~\a[120]  & ~\b[120] ;
  assign n1343 = \a[120]  & \b[120] ;
  assign n1344 = ~n1342 & ~n1343;
  assign n1345 = n1341 & ~n1344;
  assign n1346 = ~n1341 & n1344;
  assign \f[120]  = ~n1345 & ~n1346;
  assign n1348 = ~n1341 & ~n1342;
  assign n1349 = ~n1343 & ~n1348;
  assign n1350 = ~\a[121]  & ~\b[121] ;
  assign n1351 = \a[121]  & \b[121] ;
  assign n1352 = ~n1350 & ~n1351;
  assign n1353 = n1349 & ~n1352;
  assign n1354 = ~n1349 & n1352;
  assign \f[121]  = ~n1353 & ~n1354;
  assign n1356 = ~n1349 & ~n1350;
  assign n1357 = ~n1351 & ~n1356;
  assign n1358 = ~\a[122]  & ~\b[122] ;
  assign n1359 = \a[122]  & \b[122] ;
  assign n1360 = ~n1358 & ~n1359;
  assign n1361 = n1357 & ~n1360;
  assign n1362 = ~n1357 & n1360;
  assign \f[122]  = ~n1361 & ~n1362;
  assign n1364 = ~n1357 & ~n1358;
  assign n1365 = ~n1359 & ~n1364;
  assign n1366 = ~\a[123]  & ~\b[123] ;
  assign n1367 = \a[123]  & \b[123] ;
  assign n1368 = ~n1366 & ~n1367;
  assign n1369 = n1365 & ~n1368;
  assign n1370 = ~n1365 & n1368;
  assign \f[123]  = ~n1369 & ~n1370;
  assign n1372 = ~n1365 & ~n1366;
  assign n1373 = ~n1367 & ~n1372;
  assign n1374 = ~\a[124]  & ~\b[124] ;
  assign n1375 = \a[124]  & \b[124] ;
  assign n1376 = ~n1374 & ~n1375;
  assign n1377 = n1373 & ~n1376;
  assign n1378 = ~n1373 & n1376;
  assign \f[124]  = ~n1377 & ~n1378;
  assign n1380 = ~n1373 & ~n1374;
  assign n1381 = ~n1375 & ~n1380;
  assign n1382 = ~\a[125]  & ~\b[125] ;
  assign n1383 = \a[125]  & \b[125] ;
  assign n1384 = ~n1382 & ~n1383;
  assign n1385 = n1381 & ~n1384;
  assign n1386 = ~n1381 & n1384;
  assign \f[125]  = ~n1385 & ~n1386;
  assign n1388 = ~n1381 & ~n1382;
  assign n1389 = ~n1383 & ~n1388;
  assign n1390 = ~\a[126]  & ~\b[126] ;
  assign n1391 = \a[126]  & \b[126] ;
  assign n1392 = ~n1390 & ~n1391;
  assign n1393 = n1389 & ~n1392;
  assign n1394 = ~n1389 & n1392;
  assign \f[126]  = ~n1393 & ~n1394;
  assign n1396 = ~n1389 & ~n1390;
  assign n1397 = ~n1391 & ~n1396;
  assign n1398 = ~\a[127]  & ~\b[127] ;
  assign n1399 = \a[127]  & \b[127] ;
  assign n1400 = ~n1398 & ~n1399;
  assign n1401 = n1397 & ~n1400;
  assign n1402 = ~n1397 & n1400;
  assign \f[127]  = ~n1401 & ~n1402;
  assign n1404 = ~n1397 & ~n1398;
  assign cOut = n1399 | n1404;
endmodule